-- Version: 9.1 SP5 9.1.5.1
-- VHDL Black Box file 
-- 

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity roc_block is
   port( 
       RST : in std_logic;
       BCO_CLK : in std_logic;
       CLK : in std_logic;
       CLK90 : in std_logic;
       OUT_CLK : in std_logic;
       LATCH : in std_logic;
       SEND_DATA_0 : in std_logic;
       SEND_DATA_1 : in std_logic;
       DATA_IN_0 : in std_logic_vector(71 downto 0);
       DATA_IN_1 : in std_logic_vector(103 downto 0);
       SHIFT_IN : in std_logic;
       SHIFT_EN : in std_logic;
       SHIFT_OUT : out std_logic;
       LSB : out std_logic_vector(7 downto 0);
       MSB : out std_logic_vector(7 downto 0);
       DATA_OUT_0 : out std_logic_vector(31 downto 0);
       DATA_OUT_1 : out std_logic_vector(31 downto 0);
       DATA_OUT_2 : out std_logic_vector(31 downto 0);
       DATA_OUT_3 : out std_logic_vector(31 downto 0);
       TEST_OUT : out std_logic_vector(7 downto 0)
   );
end roc_block;
architecture DEF_ARCH of roc_block is 

   attribute syn_black_box : boolean;
   attribute syn_black_box of DEF_ARCH : architecture is true;
   attribute syn_tsu0: string;
   attribute syn_tsu0 of DEF_ARCH : architecture is " DATA_IN_0[0]->CLK = 1.335";
   attribute syn_tsu1: string;
   attribute syn_tsu1 of DEF_ARCH : architecture is " DATA_IN_0[0]->CLK90 = 1.33";
   attribute syn_tsu2: string;
   attribute syn_tsu2 of DEF_ARCH : architecture is " DATA_IN_0[10]->CLK = 1.335";
   attribute syn_tsu3: string;
   attribute syn_tsu3 of DEF_ARCH : architecture is " DATA_IN_0[10]->CLK90 = 1.33";
   attribute syn_tsu4: string;
   attribute syn_tsu4 of DEF_ARCH : architecture is " DATA_IN_0[11]->CLK = 1.335";
   attribute syn_tsu5: string;
   attribute syn_tsu5 of DEF_ARCH : architecture is " DATA_IN_0[11]->CLK90 = 1.33";
   attribute syn_tsu6: string;
   attribute syn_tsu6 of DEF_ARCH : architecture is " DATA_IN_0[12]->CLK = 1.335";
   attribute syn_tsu7: string;
   attribute syn_tsu7 of DEF_ARCH : architecture is " DATA_IN_0[12]->CLK90 = 1.33";
   attribute syn_tsu8: string;
   attribute syn_tsu8 of DEF_ARCH : architecture is " DATA_IN_0[13]->CLK = 1.335";
   attribute syn_tsu9: string;
   attribute syn_tsu9 of DEF_ARCH : architecture is " DATA_IN_0[13]->CLK90 = 1.33";
   attribute syn_tsu10: string;
   attribute syn_tsu10 of DEF_ARCH : architecture is " DATA_IN_0[14]->CLK = 1.335";
   attribute syn_tsu11: string;
   attribute syn_tsu11 of DEF_ARCH : architecture is " DATA_IN_0[14]->CLK90 = 1.33";
   attribute syn_tsu12: string;
   attribute syn_tsu12 of DEF_ARCH : architecture is " DATA_IN_0[15]->CLK = 1.335";
   attribute syn_tsu13: string;
   attribute syn_tsu13 of DEF_ARCH : architecture is " DATA_IN_0[15]->CLK90 = 1.33";
   attribute syn_tsu14: string;
   attribute syn_tsu14 of DEF_ARCH : architecture is " DATA_IN_0[16]->CLK = 1.335";
   attribute syn_tsu15: string;
   attribute syn_tsu15 of DEF_ARCH : architecture is " DATA_IN_0[16]->CLK90 = 1.33";
   attribute syn_tsu16: string;
   attribute syn_tsu16 of DEF_ARCH : architecture is " DATA_IN_0[17]->CLK = 1.335";
   attribute syn_tsu17: string;
   attribute syn_tsu17 of DEF_ARCH : architecture is " DATA_IN_0[17]->CLK90 = 1.33";
   attribute syn_tsu18: string;
   attribute syn_tsu18 of DEF_ARCH : architecture is " DATA_IN_0[18]->CLK = 1.335";
   attribute syn_tsu19: string;
   attribute syn_tsu19 of DEF_ARCH : architecture is " DATA_IN_0[18]->CLK90 = 1.33";
   attribute syn_tsu20: string;
   attribute syn_tsu20 of DEF_ARCH : architecture is " DATA_IN_0[19]->CLK = 1.335";
   attribute syn_tsu21: string;
   attribute syn_tsu21 of DEF_ARCH : architecture is " DATA_IN_0[19]->CLK90 = 1.33";
   attribute syn_tsu22: string;
   attribute syn_tsu22 of DEF_ARCH : architecture is " DATA_IN_0[1]->CLK = 1.335";
   attribute syn_tsu23: string;
   attribute syn_tsu23 of DEF_ARCH : architecture is " DATA_IN_0[1]->CLK90 = 1.33";
   attribute syn_tsu24: string;
   attribute syn_tsu24 of DEF_ARCH : architecture is " DATA_IN_0[20]->CLK = 1.335";
   attribute syn_tsu25: string;
   attribute syn_tsu25 of DEF_ARCH : architecture is " DATA_IN_0[20]->CLK90 = 1.33";
   attribute syn_tsu26: string;
   attribute syn_tsu26 of DEF_ARCH : architecture is " DATA_IN_0[21]->CLK = 1.335";
   attribute syn_tsu27: string;
   attribute syn_tsu27 of DEF_ARCH : architecture is " DATA_IN_0[21]->CLK90 = 1.33";
   attribute syn_tsu28: string;
   attribute syn_tsu28 of DEF_ARCH : architecture is " DATA_IN_0[22]->CLK = 1.335";
   attribute syn_tsu29: string;
   attribute syn_tsu29 of DEF_ARCH : architecture is " DATA_IN_0[22]->CLK90 = 1.33";
   attribute syn_tsu30: string;
   attribute syn_tsu30 of DEF_ARCH : architecture is " DATA_IN_0[23]->CLK = 1.335";
   attribute syn_tsu31: string;
   attribute syn_tsu31 of DEF_ARCH : architecture is " DATA_IN_0[23]->CLK90 = 1.33";
   attribute syn_tsu32: string;
   attribute syn_tsu32 of DEF_ARCH : architecture is " DATA_IN_0[24]->CLK = 1.335";
   attribute syn_tsu33: string;
   attribute syn_tsu33 of DEF_ARCH : architecture is " DATA_IN_0[24]->CLK90 = 1.33";
   attribute syn_tsu34: string;
   attribute syn_tsu34 of DEF_ARCH : architecture is " DATA_IN_0[25]->CLK = 1.335";
   attribute syn_tsu35: string;
   attribute syn_tsu35 of DEF_ARCH : architecture is " DATA_IN_0[25]->CLK90 = 1.33";
   attribute syn_tsu36: string;
   attribute syn_tsu36 of DEF_ARCH : architecture is " DATA_IN_0[26]->CLK = 1.335";
   attribute syn_tsu37: string;
   attribute syn_tsu37 of DEF_ARCH : architecture is " DATA_IN_0[26]->CLK90 = 1.33";
   attribute syn_tsu38: string;
   attribute syn_tsu38 of DEF_ARCH : architecture is " DATA_IN_0[27]->CLK = 1.335";
   attribute syn_tsu39: string;
   attribute syn_tsu39 of DEF_ARCH : architecture is " DATA_IN_0[27]->CLK90 = 1.33";
   attribute syn_tsu40: string;
   attribute syn_tsu40 of DEF_ARCH : architecture is " DATA_IN_0[28]->CLK = 1.335";
   attribute syn_tsu41: string;
   attribute syn_tsu41 of DEF_ARCH : architecture is " DATA_IN_0[28]->CLK90 = 1.33";
   attribute syn_tsu42: string;
   attribute syn_tsu42 of DEF_ARCH : architecture is " DATA_IN_0[29]->CLK = 1.335";
   attribute syn_tsu43: string;
   attribute syn_tsu43 of DEF_ARCH : architecture is " DATA_IN_0[29]->CLK90 = 1.33";
   attribute syn_tsu44: string;
   attribute syn_tsu44 of DEF_ARCH : architecture is " DATA_IN_0[2]->CLK = 1.335";
   attribute syn_tsu45: string;
   attribute syn_tsu45 of DEF_ARCH : architecture is " DATA_IN_0[2]->CLK90 = 1.33";
   attribute syn_tsu46: string;
   attribute syn_tsu46 of DEF_ARCH : architecture is " DATA_IN_0[30]->CLK = 1.335";
   attribute syn_tsu47: string;
   attribute syn_tsu47 of DEF_ARCH : architecture is " DATA_IN_0[30]->CLK90 = 1.33";
   attribute syn_tsu48: string;
   attribute syn_tsu48 of DEF_ARCH : architecture is " DATA_IN_0[31]->CLK = 1.335";
   attribute syn_tsu49: string;
   attribute syn_tsu49 of DEF_ARCH : architecture is " DATA_IN_0[31]->CLK90 = 1.33";
   attribute syn_tsu50: string;
   attribute syn_tsu50 of DEF_ARCH : architecture is " DATA_IN_0[32]->CLK = 1.335";
   attribute syn_tsu51: string;
   attribute syn_tsu51 of DEF_ARCH : architecture is " DATA_IN_0[32]->CLK90 = 1.33";
   attribute syn_tsu52: string;
   attribute syn_tsu52 of DEF_ARCH : architecture is " DATA_IN_0[33]->CLK = 1.335";
   attribute syn_tsu53: string;
   attribute syn_tsu53 of DEF_ARCH : architecture is " DATA_IN_0[33]->CLK90 = 1.33";
   attribute syn_tsu54: string;
   attribute syn_tsu54 of DEF_ARCH : architecture is " DATA_IN_0[34]->CLK = 1.335";
   attribute syn_tsu55: string;
   attribute syn_tsu55 of DEF_ARCH : architecture is " DATA_IN_0[34]->CLK90 = 1.33";
   attribute syn_tsu56: string;
   attribute syn_tsu56 of DEF_ARCH : architecture is " DATA_IN_0[35]->CLK = 1.335";
   attribute syn_tsu57: string;
   attribute syn_tsu57 of DEF_ARCH : architecture is " DATA_IN_0[35]->CLK90 = 1.33";
   attribute syn_tsu58: string;
   attribute syn_tsu58 of DEF_ARCH : architecture is " DATA_IN_0[36]->CLK = 1.335";
   attribute syn_tsu59: string;
   attribute syn_tsu59 of DEF_ARCH : architecture is " DATA_IN_0[36]->CLK90 = 1.33";
   attribute syn_tsu60: string;
   attribute syn_tsu60 of DEF_ARCH : architecture is " DATA_IN_0[37]->CLK = 1.335";
   attribute syn_tsu61: string;
   attribute syn_tsu61 of DEF_ARCH : architecture is " DATA_IN_0[37]->CLK90 = 1.33";
   attribute syn_tsu62: string;
   attribute syn_tsu62 of DEF_ARCH : architecture is " DATA_IN_0[38]->CLK = 1.335";
   attribute syn_tsu63: string;
   attribute syn_tsu63 of DEF_ARCH : architecture is " DATA_IN_0[38]->CLK90 = 1.33";
   attribute syn_tsu64: string;
   attribute syn_tsu64 of DEF_ARCH : architecture is " DATA_IN_0[39]->CLK = 1.335";
   attribute syn_tsu65: string;
   attribute syn_tsu65 of DEF_ARCH : architecture is " DATA_IN_0[39]->CLK90 = 1.33";
   attribute syn_tsu66: string;
   attribute syn_tsu66 of DEF_ARCH : architecture is " DATA_IN_0[3]->CLK = 1.335";
   attribute syn_tsu67: string;
   attribute syn_tsu67 of DEF_ARCH : architecture is " DATA_IN_0[3]->CLK90 = 1.33";
   attribute syn_tsu68: string;
   attribute syn_tsu68 of DEF_ARCH : architecture is " DATA_IN_0[40]->CLK = 1.335";
   attribute syn_tsu69: string;
   attribute syn_tsu69 of DEF_ARCH : architecture is " DATA_IN_0[40]->CLK90 = 1.33";
   attribute syn_tsu70: string;
   attribute syn_tsu70 of DEF_ARCH : architecture is " DATA_IN_0[41]->CLK = 1.335";
   attribute syn_tsu71: string;
   attribute syn_tsu71 of DEF_ARCH : architecture is " DATA_IN_0[41]->CLK90 = 1.33";
   attribute syn_tsu72: string;
   attribute syn_tsu72 of DEF_ARCH : architecture is " DATA_IN_0[42]->CLK = 1.335";
   attribute syn_tsu73: string;
   attribute syn_tsu73 of DEF_ARCH : architecture is " DATA_IN_0[42]->CLK90 = 1.33";
   attribute syn_tsu74: string;
   attribute syn_tsu74 of DEF_ARCH : architecture is " DATA_IN_0[43]->CLK = 1.335";
   attribute syn_tsu75: string;
   attribute syn_tsu75 of DEF_ARCH : architecture is " DATA_IN_0[43]->CLK90 = 1.33";
   attribute syn_tsu76: string;
   attribute syn_tsu76 of DEF_ARCH : architecture is " DATA_IN_0[44]->CLK = 1.335";
   attribute syn_tsu77: string;
   attribute syn_tsu77 of DEF_ARCH : architecture is " DATA_IN_0[44]->CLK90 = 1.33";
   attribute syn_tsu78: string;
   attribute syn_tsu78 of DEF_ARCH : architecture is " DATA_IN_0[45]->CLK = 1.335";
   attribute syn_tsu79: string;
   attribute syn_tsu79 of DEF_ARCH : architecture is " DATA_IN_0[45]->CLK90 = 1.33";
   attribute syn_tsu80: string;
   attribute syn_tsu80 of DEF_ARCH : architecture is " DATA_IN_0[46]->CLK = 1.335";
   attribute syn_tsu81: string;
   attribute syn_tsu81 of DEF_ARCH : architecture is " DATA_IN_0[46]->CLK90 = 1.33";
   attribute syn_tsu82: string;
   attribute syn_tsu82 of DEF_ARCH : architecture is " DATA_IN_0[47]->CLK = 1.335";
   attribute syn_tsu83: string;
   attribute syn_tsu83 of DEF_ARCH : architecture is " DATA_IN_0[47]->CLK90 = 1.33";
   attribute syn_tsu84: string;
   attribute syn_tsu84 of DEF_ARCH : architecture is " DATA_IN_0[48]->CLK = 1.335";
   attribute syn_tsu85: string;
   attribute syn_tsu85 of DEF_ARCH : architecture is " DATA_IN_0[48]->CLK90 = 1.33";
   attribute syn_tsu86: string;
   attribute syn_tsu86 of DEF_ARCH : architecture is " DATA_IN_0[49]->CLK = 1.335";
   attribute syn_tsu87: string;
   attribute syn_tsu87 of DEF_ARCH : architecture is " DATA_IN_0[49]->CLK90 = 1.33";
   attribute syn_tsu88: string;
   attribute syn_tsu88 of DEF_ARCH : architecture is " DATA_IN_0[4]->CLK = 1.335";
   attribute syn_tsu89: string;
   attribute syn_tsu89 of DEF_ARCH : architecture is " DATA_IN_0[4]->CLK90 = 1.33";
   attribute syn_tsu90: string;
   attribute syn_tsu90 of DEF_ARCH : architecture is " DATA_IN_0[50]->CLK = 1.335";
   attribute syn_tsu91: string;
   attribute syn_tsu91 of DEF_ARCH : architecture is " DATA_IN_0[50]->CLK90 = 1.33";
   attribute syn_tsu92: string;
   attribute syn_tsu92 of DEF_ARCH : architecture is " DATA_IN_0[51]->CLK = 1.335";
   attribute syn_tsu93: string;
   attribute syn_tsu93 of DEF_ARCH : architecture is " DATA_IN_0[51]->CLK90 = 1.33";
   attribute syn_tsu94: string;
   attribute syn_tsu94 of DEF_ARCH : architecture is " DATA_IN_0[52]->CLK = 1.335";
   attribute syn_tsu95: string;
   attribute syn_tsu95 of DEF_ARCH : architecture is " DATA_IN_0[52]->CLK90 = 1.33";
   attribute syn_tsu96: string;
   attribute syn_tsu96 of DEF_ARCH : architecture is " DATA_IN_0[53]->CLK = 1.335";
   attribute syn_tsu97: string;
   attribute syn_tsu97 of DEF_ARCH : architecture is " DATA_IN_0[53]->CLK90 = 1.33";
   attribute syn_tsu98: string;
   attribute syn_tsu98 of DEF_ARCH : architecture is " DATA_IN_0[54]->CLK = 1.335";
   attribute syn_tsu99: string;
   attribute syn_tsu99 of DEF_ARCH : architecture is " DATA_IN_0[54]->CLK90 = 1.33";
   attribute syn_tsu100: string;
   attribute syn_tsu100 of DEF_ARCH : architecture is " DATA_IN_0[55]->CLK = 1.335";
   attribute syn_tsu101: string;
   attribute syn_tsu101 of DEF_ARCH : architecture is " DATA_IN_0[55]->CLK90 = 1.33";
   attribute syn_tsu102: string;
   attribute syn_tsu102 of DEF_ARCH : architecture is " DATA_IN_0[56]->CLK = 1.335";
   attribute syn_tsu103: string;
   attribute syn_tsu103 of DEF_ARCH : architecture is " DATA_IN_0[56]->CLK90 = 1.33";
   attribute syn_tsu104: string;
   attribute syn_tsu104 of DEF_ARCH : architecture is " DATA_IN_0[57]->CLK = 1.335";
   attribute syn_tsu105: string;
   attribute syn_tsu105 of DEF_ARCH : architecture is " DATA_IN_0[57]->CLK90 = 1.33";
   attribute syn_tsu106: string;
   attribute syn_tsu106 of DEF_ARCH : architecture is " DATA_IN_0[58]->CLK = 1.335";
   attribute syn_tsu107: string;
   attribute syn_tsu107 of DEF_ARCH : architecture is " DATA_IN_0[58]->CLK90 = 1.33";
   attribute syn_tsu108: string;
   attribute syn_tsu108 of DEF_ARCH : architecture is " DATA_IN_0[59]->CLK = 1.335";
   attribute syn_tsu109: string;
   attribute syn_tsu109 of DEF_ARCH : architecture is " DATA_IN_0[59]->CLK90 = 1.33";
   attribute syn_tsu110: string;
   attribute syn_tsu110 of DEF_ARCH : architecture is " DATA_IN_0[5]->CLK = 1.335";
   attribute syn_tsu111: string;
   attribute syn_tsu111 of DEF_ARCH : architecture is " DATA_IN_0[5]->CLK90 = 1.33";
   attribute syn_tsu112: string;
   attribute syn_tsu112 of DEF_ARCH : architecture is " DATA_IN_0[60]->CLK = 1.335";
   attribute syn_tsu113: string;
   attribute syn_tsu113 of DEF_ARCH : architecture is " DATA_IN_0[60]->CLK90 = 1.33";
   attribute syn_tsu114: string;
   attribute syn_tsu114 of DEF_ARCH : architecture is " DATA_IN_0[61]->CLK = 1.335";
   attribute syn_tsu115: string;
   attribute syn_tsu115 of DEF_ARCH : architecture is " DATA_IN_0[61]->CLK90 = 1.33";
   attribute syn_tsu116: string;
   attribute syn_tsu116 of DEF_ARCH : architecture is " DATA_IN_0[62]->CLK = 1.335";
   attribute syn_tsu117: string;
   attribute syn_tsu117 of DEF_ARCH : architecture is " DATA_IN_0[62]->CLK90 = 1.33";
   attribute syn_tsu118: string;
   attribute syn_tsu118 of DEF_ARCH : architecture is " DATA_IN_0[63]->CLK = 1.335";
   attribute syn_tsu119: string;
   attribute syn_tsu119 of DEF_ARCH : architecture is " DATA_IN_0[63]->CLK90 = 1.33";
   attribute syn_tsu120: string;
   attribute syn_tsu120 of DEF_ARCH : architecture is " DATA_IN_0[64]->CLK = 1.335";
   attribute syn_tsu121: string;
   attribute syn_tsu121 of DEF_ARCH : architecture is " DATA_IN_0[64]->CLK90 = 1.33";
   attribute syn_tsu122: string;
   attribute syn_tsu122 of DEF_ARCH : architecture is " DATA_IN_0[65]->CLK = 1.335";
   attribute syn_tsu123: string;
   attribute syn_tsu123 of DEF_ARCH : architecture is " DATA_IN_0[65]->CLK90 = 1.33";
   attribute syn_tsu124: string;
   attribute syn_tsu124 of DEF_ARCH : architecture is " DATA_IN_0[66]->CLK = 1.335";
   attribute syn_tsu125: string;
   attribute syn_tsu125 of DEF_ARCH : architecture is " DATA_IN_0[66]->CLK90 = 1.33";
   attribute syn_tsu126: string;
   attribute syn_tsu126 of DEF_ARCH : architecture is " DATA_IN_0[67]->CLK = 1.335";
   attribute syn_tsu127: string;
   attribute syn_tsu127 of DEF_ARCH : architecture is " DATA_IN_0[67]->CLK90 = 1.33";
   attribute syn_tsu128: string;
   attribute syn_tsu128 of DEF_ARCH : architecture is " DATA_IN_0[68]->CLK = 1.335";
   attribute syn_tsu129: string;
   attribute syn_tsu129 of DEF_ARCH : architecture is " DATA_IN_0[68]->CLK90 = 1.33";
   attribute syn_tsu130: string;
   attribute syn_tsu130 of DEF_ARCH : architecture is " DATA_IN_0[69]->CLK = 1.335";
   attribute syn_tsu131: string;
   attribute syn_tsu131 of DEF_ARCH : architecture is " DATA_IN_0[69]->CLK90 = 1.33";
   attribute syn_tsu132: string;
   attribute syn_tsu132 of DEF_ARCH : architecture is " DATA_IN_0[6]->CLK = 1.335";
   attribute syn_tsu133: string;
   attribute syn_tsu133 of DEF_ARCH : architecture is " DATA_IN_0[6]->CLK90 = 1.33";
   attribute syn_tsu134: string;
   attribute syn_tsu134 of DEF_ARCH : architecture is " DATA_IN_0[70]->CLK = 1.335";
   attribute syn_tsu135: string;
   attribute syn_tsu135 of DEF_ARCH : architecture is " DATA_IN_0[70]->CLK90 = 1.33";
   attribute syn_tsu136: string;
   attribute syn_tsu136 of DEF_ARCH : architecture is " DATA_IN_0[71]->CLK = 1.335";
   attribute syn_tsu137: string;
   attribute syn_tsu137 of DEF_ARCH : architecture is " DATA_IN_0[71]->CLK90 = 1.33";
   attribute syn_tsu138: string;
   attribute syn_tsu138 of DEF_ARCH : architecture is " DATA_IN_0[7]->CLK = 1.335";
   attribute syn_tsu139: string;
   attribute syn_tsu139 of DEF_ARCH : architecture is " DATA_IN_0[7]->CLK90 = 1.33";
   attribute syn_tsu140: string;
   attribute syn_tsu140 of DEF_ARCH : architecture is " DATA_IN_0[8]->CLK = 1.335";
   attribute syn_tsu141: string;
   attribute syn_tsu141 of DEF_ARCH : architecture is " DATA_IN_0[8]->CLK90 = 1.33";
   attribute syn_tsu142: string;
   attribute syn_tsu142 of DEF_ARCH : architecture is " DATA_IN_0[9]->CLK = 1.335";
   attribute syn_tsu143: string;
   attribute syn_tsu143 of DEF_ARCH : architecture is " DATA_IN_0[9]->CLK90 = 1.33";
   attribute syn_tsu144: string;
   attribute syn_tsu144 of DEF_ARCH : architecture is " DATA_IN_1[0]->CLK = 1.335";
   attribute syn_tsu145: string;
   attribute syn_tsu145 of DEF_ARCH : architecture is " DATA_IN_1[0]->CLK90 = 1.33";
   attribute syn_tsu146: string;
   attribute syn_tsu146 of DEF_ARCH : architecture is " DATA_IN_1[100]->CLK = 1.335";
   attribute syn_tsu147: string;
   attribute syn_tsu147 of DEF_ARCH : architecture is " DATA_IN_1[100]->CLK90 = 1.33";
   attribute syn_tsu148: string;
   attribute syn_tsu148 of DEF_ARCH : architecture is " DATA_IN_1[101]->CLK = 1.335";
   attribute syn_tsu149: string;
   attribute syn_tsu149 of DEF_ARCH : architecture is " DATA_IN_1[101]->CLK90 = 1.33";
   attribute syn_tsu150: string;
   attribute syn_tsu150 of DEF_ARCH : architecture is " DATA_IN_1[102]->CLK = 1.335";
   attribute syn_tsu151: string;
   attribute syn_tsu151 of DEF_ARCH : architecture is " DATA_IN_1[102]->CLK90 = 1.33";
   attribute syn_tsu152: string;
   attribute syn_tsu152 of DEF_ARCH : architecture is " DATA_IN_1[103]->CLK = 1.335";
   attribute syn_tsu153: string;
   attribute syn_tsu153 of DEF_ARCH : architecture is " DATA_IN_1[103]->CLK90 = 1.33";
   attribute syn_tsu154: string;
   attribute syn_tsu154 of DEF_ARCH : architecture is " DATA_IN_1[10]->CLK = 1.335";
   attribute syn_tsu155: string;
   attribute syn_tsu155 of DEF_ARCH : architecture is " DATA_IN_1[10]->CLK90 = 1.33";
   attribute syn_tsu156: string;
   attribute syn_tsu156 of DEF_ARCH : architecture is " DATA_IN_1[11]->CLK = 1.335";
   attribute syn_tsu157: string;
   attribute syn_tsu157 of DEF_ARCH : architecture is " DATA_IN_1[11]->CLK90 = 1.33";
   attribute syn_tsu158: string;
   attribute syn_tsu158 of DEF_ARCH : architecture is " DATA_IN_1[12]->CLK = 1.335";
   attribute syn_tsu159: string;
   attribute syn_tsu159 of DEF_ARCH : architecture is " DATA_IN_1[12]->CLK90 = 1.33";
   attribute syn_tsu160: string;
   attribute syn_tsu160 of DEF_ARCH : architecture is " DATA_IN_1[13]->CLK = 1.335";
   attribute syn_tsu161: string;
   attribute syn_tsu161 of DEF_ARCH : architecture is " DATA_IN_1[13]->CLK90 = 1.33";
   attribute syn_tsu162: string;
   attribute syn_tsu162 of DEF_ARCH : architecture is " DATA_IN_1[14]->CLK = 1.335";
   attribute syn_tsu163: string;
   attribute syn_tsu163 of DEF_ARCH : architecture is " DATA_IN_1[14]->CLK90 = 1.33";
   attribute syn_tsu164: string;
   attribute syn_tsu164 of DEF_ARCH : architecture is " DATA_IN_1[15]->CLK = 1.335";
   attribute syn_tsu165: string;
   attribute syn_tsu165 of DEF_ARCH : architecture is " DATA_IN_1[15]->CLK90 = 1.33";
   attribute syn_tsu166: string;
   attribute syn_tsu166 of DEF_ARCH : architecture is " DATA_IN_1[16]->CLK = 1.335";
   attribute syn_tsu167: string;
   attribute syn_tsu167 of DEF_ARCH : architecture is " DATA_IN_1[16]->CLK90 = 1.33";
   attribute syn_tsu168: string;
   attribute syn_tsu168 of DEF_ARCH : architecture is " DATA_IN_1[17]->CLK = 1.335";
   attribute syn_tsu169: string;
   attribute syn_tsu169 of DEF_ARCH : architecture is " DATA_IN_1[17]->CLK90 = 1.33";
   attribute syn_tsu170: string;
   attribute syn_tsu170 of DEF_ARCH : architecture is " DATA_IN_1[18]->CLK = 1.335";
   attribute syn_tsu171: string;
   attribute syn_tsu171 of DEF_ARCH : architecture is " DATA_IN_1[18]->CLK90 = 1.33";
   attribute syn_tsu172: string;
   attribute syn_tsu172 of DEF_ARCH : architecture is " DATA_IN_1[19]->CLK = 1.335";
   attribute syn_tsu173: string;
   attribute syn_tsu173 of DEF_ARCH : architecture is " DATA_IN_1[19]->CLK90 = 1.33";
   attribute syn_tsu174: string;
   attribute syn_tsu174 of DEF_ARCH : architecture is " DATA_IN_1[1]->CLK = 1.335";
   attribute syn_tsu175: string;
   attribute syn_tsu175 of DEF_ARCH : architecture is " DATA_IN_1[1]->CLK90 = 1.33";
   attribute syn_tsu176: string;
   attribute syn_tsu176 of DEF_ARCH : architecture is " DATA_IN_1[20]->CLK = 1.335";
   attribute syn_tsu177: string;
   attribute syn_tsu177 of DEF_ARCH : architecture is " DATA_IN_1[20]->CLK90 = 1.33";
   attribute syn_tsu178: string;
   attribute syn_tsu178 of DEF_ARCH : architecture is " DATA_IN_1[21]->CLK = 1.335";
   attribute syn_tsu179: string;
   attribute syn_tsu179 of DEF_ARCH : architecture is " DATA_IN_1[21]->CLK90 = 1.33";
   attribute syn_tsu180: string;
   attribute syn_tsu180 of DEF_ARCH : architecture is " DATA_IN_1[22]->CLK = 1.335";
   attribute syn_tsu181: string;
   attribute syn_tsu181 of DEF_ARCH : architecture is " DATA_IN_1[22]->CLK90 = 1.33";
   attribute syn_tsu182: string;
   attribute syn_tsu182 of DEF_ARCH : architecture is " DATA_IN_1[23]->CLK = 1.335";
   attribute syn_tsu183: string;
   attribute syn_tsu183 of DEF_ARCH : architecture is " DATA_IN_1[23]->CLK90 = 1.33";
   attribute syn_tsu184: string;
   attribute syn_tsu184 of DEF_ARCH : architecture is " DATA_IN_1[24]->CLK = 1.335";
   attribute syn_tsu185: string;
   attribute syn_tsu185 of DEF_ARCH : architecture is " DATA_IN_1[24]->CLK90 = 1.33";
   attribute syn_tsu186: string;
   attribute syn_tsu186 of DEF_ARCH : architecture is " DATA_IN_1[25]->CLK = 1.335";
   attribute syn_tsu187: string;
   attribute syn_tsu187 of DEF_ARCH : architecture is " DATA_IN_1[25]->CLK90 = 1.33";
   attribute syn_tsu188: string;
   attribute syn_tsu188 of DEF_ARCH : architecture is " DATA_IN_1[26]->CLK = 1.335";
   attribute syn_tsu189: string;
   attribute syn_tsu189 of DEF_ARCH : architecture is " DATA_IN_1[26]->CLK90 = 1.33";
   attribute syn_tsu190: string;
   attribute syn_tsu190 of DEF_ARCH : architecture is " DATA_IN_1[27]->CLK = 1.335";
   attribute syn_tsu191: string;
   attribute syn_tsu191 of DEF_ARCH : architecture is " DATA_IN_1[27]->CLK90 = 1.33";
   attribute syn_tsu192: string;
   attribute syn_tsu192 of DEF_ARCH : architecture is " DATA_IN_1[28]->CLK = 1.335";
   attribute syn_tsu193: string;
   attribute syn_tsu193 of DEF_ARCH : architecture is " DATA_IN_1[28]->CLK90 = 1.33";
   attribute syn_tsu194: string;
   attribute syn_tsu194 of DEF_ARCH : architecture is " DATA_IN_1[29]->CLK = 1.335";
   attribute syn_tsu195: string;
   attribute syn_tsu195 of DEF_ARCH : architecture is " DATA_IN_1[29]->CLK90 = 1.33";
   attribute syn_tsu196: string;
   attribute syn_tsu196 of DEF_ARCH : architecture is " DATA_IN_1[2]->CLK = 1.335";
   attribute syn_tsu197: string;
   attribute syn_tsu197 of DEF_ARCH : architecture is " DATA_IN_1[2]->CLK90 = 1.33";
   attribute syn_tsu198: string;
   attribute syn_tsu198 of DEF_ARCH : architecture is " DATA_IN_1[30]->CLK = 1.335";
   attribute syn_tsu199: string;
   attribute syn_tsu199 of DEF_ARCH : architecture is " DATA_IN_1[30]->CLK90 = 1.33";
   attribute syn_tsu200: string;
   attribute syn_tsu200 of DEF_ARCH : architecture is " DATA_IN_1[31]->CLK = 1.335";
   attribute syn_tsu201: string;
   attribute syn_tsu201 of DEF_ARCH : architecture is " DATA_IN_1[31]->CLK90 = 1.33";
   attribute syn_tsu202: string;
   attribute syn_tsu202 of DEF_ARCH : architecture is " DATA_IN_1[32]->CLK = 1.335";
   attribute syn_tsu203: string;
   attribute syn_tsu203 of DEF_ARCH : architecture is " DATA_IN_1[32]->CLK90 = 1.33";
   attribute syn_tsu204: string;
   attribute syn_tsu204 of DEF_ARCH : architecture is " DATA_IN_1[33]->CLK = 1.335";
   attribute syn_tsu205: string;
   attribute syn_tsu205 of DEF_ARCH : architecture is " DATA_IN_1[33]->CLK90 = 1.33";
   attribute syn_tsu206: string;
   attribute syn_tsu206 of DEF_ARCH : architecture is " DATA_IN_1[34]->CLK = 1.335";
   attribute syn_tsu207: string;
   attribute syn_tsu207 of DEF_ARCH : architecture is " DATA_IN_1[34]->CLK90 = 1.33";
   attribute syn_tsu208: string;
   attribute syn_tsu208 of DEF_ARCH : architecture is " DATA_IN_1[35]->CLK = 1.335";
   attribute syn_tsu209: string;
   attribute syn_tsu209 of DEF_ARCH : architecture is " DATA_IN_1[35]->CLK90 = 1.33";
   attribute syn_tsu210: string;
   attribute syn_tsu210 of DEF_ARCH : architecture is " DATA_IN_1[36]->CLK = 1.335";
   attribute syn_tsu211: string;
   attribute syn_tsu211 of DEF_ARCH : architecture is " DATA_IN_1[36]->CLK90 = 1.33";
   attribute syn_tsu212: string;
   attribute syn_tsu212 of DEF_ARCH : architecture is " DATA_IN_1[37]->CLK = 1.335";
   attribute syn_tsu213: string;
   attribute syn_tsu213 of DEF_ARCH : architecture is " DATA_IN_1[37]->CLK90 = 1.33";
   attribute syn_tsu214: string;
   attribute syn_tsu214 of DEF_ARCH : architecture is " DATA_IN_1[38]->CLK = 1.335";
   attribute syn_tsu215: string;
   attribute syn_tsu215 of DEF_ARCH : architecture is " DATA_IN_1[38]->CLK90 = 1.33";
   attribute syn_tsu216: string;
   attribute syn_tsu216 of DEF_ARCH : architecture is " DATA_IN_1[39]->CLK = 1.335";
   attribute syn_tsu217: string;
   attribute syn_tsu217 of DEF_ARCH : architecture is " DATA_IN_1[39]->CLK90 = 1.33";
   attribute syn_tsu218: string;
   attribute syn_tsu218 of DEF_ARCH : architecture is " DATA_IN_1[3]->CLK = 1.335";
   attribute syn_tsu219: string;
   attribute syn_tsu219 of DEF_ARCH : architecture is " DATA_IN_1[3]->CLK90 = 1.33";
   attribute syn_tsu220: string;
   attribute syn_tsu220 of DEF_ARCH : architecture is " DATA_IN_1[40]->CLK = 1.335";
   attribute syn_tsu221: string;
   attribute syn_tsu221 of DEF_ARCH : architecture is " DATA_IN_1[40]->CLK90 = 1.33";
   attribute syn_tsu222: string;
   attribute syn_tsu222 of DEF_ARCH : architecture is " DATA_IN_1[41]->CLK = 1.335";
   attribute syn_tsu223: string;
   attribute syn_tsu223 of DEF_ARCH : architecture is " DATA_IN_1[41]->CLK90 = 1.33";
   attribute syn_tsu224: string;
   attribute syn_tsu224 of DEF_ARCH : architecture is " DATA_IN_1[42]->CLK = 1.335";
   attribute syn_tsu225: string;
   attribute syn_tsu225 of DEF_ARCH : architecture is " DATA_IN_1[42]->CLK90 = 1.33";
   attribute syn_tsu226: string;
   attribute syn_tsu226 of DEF_ARCH : architecture is " DATA_IN_1[43]->CLK = 1.335";
   attribute syn_tsu227: string;
   attribute syn_tsu227 of DEF_ARCH : architecture is " DATA_IN_1[43]->CLK90 = 1.33";
   attribute syn_tsu228: string;
   attribute syn_tsu228 of DEF_ARCH : architecture is " DATA_IN_1[44]->CLK = 1.335";
   attribute syn_tsu229: string;
   attribute syn_tsu229 of DEF_ARCH : architecture is " DATA_IN_1[44]->CLK90 = 1.33";
   attribute syn_tsu230: string;
   attribute syn_tsu230 of DEF_ARCH : architecture is " DATA_IN_1[45]->CLK = 1.335";
   attribute syn_tsu231: string;
   attribute syn_tsu231 of DEF_ARCH : architecture is " DATA_IN_1[45]->CLK90 = 1.33";
   attribute syn_tsu232: string;
   attribute syn_tsu232 of DEF_ARCH : architecture is " DATA_IN_1[46]->CLK = 1.335";
   attribute syn_tsu233: string;
   attribute syn_tsu233 of DEF_ARCH : architecture is " DATA_IN_1[46]->CLK90 = 1.33";
   attribute syn_tsu234: string;
   attribute syn_tsu234 of DEF_ARCH : architecture is " DATA_IN_1[47]->CLK = 1.335";
   attribute syn_tsu235: string;
   attribute syn_tsu235 of DEF_ARCH : architecture is " DATA_IN_1[47]->CLK90 = 1.33";
   attribute syn_tsu236: string;
   attribute syn_tsu236 of DEF_ARCH : architecture is " DATA_IN_1[48]->CLK = 1.335";
   attribute syn_tsu237: string;
   attribute syn_tsu237 of DEF_ARCH : architecture is " DATA_IN_1[48]->CLK90 = 1.33";
   attribute syn_tsu238: string;
   attribute syn_tsu238 of DEF_ARCH : architecture is " DATA_IN_1[49]->CLK = 1.335";
   attribute syn_tsu239: string;
   attribute syn_tsu239 of DEF_ARCH : architecture is " DATA_IN_1[49]->CLK90 = 1.33";
   attribute syn_tsu240: string;
   attribute syn_tsu240 of DEF_ARCH : architecture is " DATA_IN_1[4]->CLK = 1.335";
   attribute syn_tsu241: string;
   attribute syn_tsu241 of DEF_ARCH : architecture is " DATA_IN_1[4]->CLK90 = 1.33";
   attribute syn_tsu242: string;
   attribute syn_tsu242 of DEF_ARCH : architecture is " DATA_IN_1[50]->CLK = 1.335";
   attribute syn_tsu243: string;
   attribute syn_tsu243 of DEF_ARCH : architecture is " DATA_IN_1[50]->CLK90 = 1.33";
   attribute syn_tsu244: string;
   attribute syn_tsu244 of DEF_ARCH : architecture is " DATA_IN_1[51]->CLK = 1.335";
   attribute syn_tsu245: string;
   attribute syn_tsu245 of DEF_ARCH : architecture is " DATA_IN_1[51]->CLK90 = 1.33";
   attribute syn_tsu246: string;
   attribute syn_tsu246 of DEF_ARCH : architecture is " DATA_IN_1[52]->CLK = 1.335";
   attribute syn_tsu247: string;
   attribute syn_tsu247 of DEF_ARCH : architecture is " DATA_IN_1[52]->CLK90 = 1.33";
   attribute syn_tsu248: string;
   attribute syn_tsu248 of DEF_ARCH : architecture is " DATA_IN_1[53]->CLK = 1.335";
   attribute syn_tsu249: string;
   attribute syn_tsu249 of DEF_ARCH : architecture is " DATA_IN_1[53]->CLK90 = 1.33";
   attribute syn_tsu250: string;
   attribute syn_tsu250 of DEF_ARCH : architecture is " DATA_IN_1[54]->CLK = 1.335";
   attribute syn_tsu251: string;
   attribute syn_tsu251 of DEF_ARCH : architecture is " DATA_IN_1[54]->CLK90 = 1.33";
   attribute syn_tsu252: string;
   attribute syn_tsu252 of DEF_ARCH : architecture is " DATA_IN_1[55]->CLK = 1.335";
   attribute syn_tsu253: string;
   attribute syn_tsu253 of DEF_ARCH : architecture is " DATA_IN_1[55]->CLK90 = 1.33";
   attribute syn_tsu254: string;
   attribute syn_tsu254 of DEF_ARCH : architecture is " DATA_IN_1[56]->CLK = 1.335";
   attribute syn_tsu255: string;
   attribute syn_tsu255 of DEF_ARCH : architecture is " DATA_IN_1[56]->CLK90 = 1.33";
   attribute syn_tsu256: string;
   attribute syn_tsu256 of DEF_ARCH : architecture is " DATA_IN_1[57]->CLK = 1.335";
   attribute syn_tsu257: string;
   attribute syn_tsu257 of DEF_ARCH : architecture is " DATA_IN_1[57]->CLK90 = 1.33";
   attribute syn_tsu258: string;
   attribute syn_tsu258 of DEF_ARCH : architecture is " DATA_IN_1[58]->CLK = 1.335";
   attribute syn_tsu259: string;
   attribute syn_tsu259 of DEF_ARCH : architecture is " DATA_IN_1[58]->CLK90 = 1.33";
   attribute syn_tsu260: string;
   attribute syn_tsu260 of DEF_ARCH : architecture is " DATA_IN_1[59]->CLK = 1.335";
   attribute syn_tsu261: string;
   attribute syn_tsu261 of DEF_ARCH : architecture is " DATA_IN_1[59]->CLK90 = 1.33";
   attribute syn_tsu262: string;
   attribute syn_tsu262 of DEF_ARCH : architecture is " DATA_IN_1[5]->CLK = 1.335";
   attribute syn_tsu263: string;
   attribute syn_tsu263 of DEF_ARCH : architecture is " DATA_IN_1[5]->CLK90 = 1.33";
   attribute syn_tsu264: string;
   attribute syn_tsu264 of DEF_ARCH : architecture is " DATA_IN_1[60]->CLK = 1.335";
   attribute syn_tsu265: string;
   attribute syn_tsu265 of DEF_ARCH : architecture is " DATA_IN_1[60]->CLK90 = 1.33";
   attribute syn_tsu266: string;
   attribute syn_tsu266 of DEF_ARCH : architecture is " DATA_IN_1[61]->CLK = 1.335";
   attribute syn_tsu267: string;
   attribute syn_tsu267 of DEF_ARCH : architecture is " DATA_IN_1[61]->CLK90 = 1.33";
   attribute syn_tsu268: string;
   attribute syn_tsu268 of DEF_ARCH : architecture is " DATA_IN_1[62]->CLK = 1.335";
   attribute syn_tsu269: string;
   attribute syn_tsu269 of DEF_ARCH : architecture is " DATA_IN_1[62]->CLK90 = 1.33";
   attribute syn_tsu270: string;
   attribute syn_tsu270 of DEF_ARCH : architecture is " DATA_IN_1[63]->CLK = 1.335";
   attribute syn_tsu271: string;
   attribute syn_tsu271 of DEF_ARCH : architecture is " DATA_IN_1[63]->CLK90 = 1.33";
   attribute syn_tsu272: string;
   attribute syn_tsu272 of DEF_ARCH : architecture is " DATA_IN_1[64]->CLK = 1.335";
   attribute syn_tsu273: string;
   attribute syn_tsu273 of DEF_ARCH : architecture is " DATA_IN_1[64]->CLK90 = 1.33";
   attribute syn_tsu274: string;
   attribute syn_tsu274 of DEF_ARCH : architecture is " DATA_IN_1[65]->CLK = 1.335";
   attribute syn_tsu275: string;
   attribute syn_tsu275 of DEF_ARCH : architecture is " DATA_IN_1[65]->CLK90 = 1.33";
   attribute syn_tsu276: string;
   attribute syn_tsu276 of DEF_ARCH : architecture is " DATA_IN_1[66]->CLK = 1.335";
   attribute syn_tsu277: string;
   attribute syn_tsu277 of DEF_ARCH : architecture is " DATA_IN_1[66]->CLK90 = 1.33";
   attribute syn_tsu278: string;
   attribute syn_tsu278 of DEF_ARCH : architecture is " DATA_IN_1[67]->CLK = 1.335";
   attribute syn_tsu279: string;
   attribute syn_tsu279 of DEF_ARCH : architecture is " DATA_IN_1[67]->CLK90 = 1.33";
   attribute syn_tsu280: string;
   attribute syn_tsu280 of DEF_ARCH : architecture is " DATA_IN_1[68]->CLK = 1.335";
   attribute syn_tsu281: string;
   attribute syn_tsu281 of DEF_ARCH : architecture is " DATA_IN_1[68]->CLK90 = 1.33";
   attribute syn_tsu282: string;
   attribute syn_tsu282 of DEF_ARCH : architecture is " DATA_IN_1[69]->CLK = 1.335";
   attribute syn_tsu283: string;
   attribute syn_tsu283 of DEF_ARCH : architecture is " DATA_IN_1[69]->CLK90 = 1.33";
   attribute syn_tsu284: string;
   attribute syn_tsu284 of DEF_ARCH : architecture is " DATA_IN_1[6]->CLK = 1.335";
   attribute syn_tsu285: string;
   attribute syn_tsu285 of DEF_ARCH : architecture is " DATA_IN_1[6]->CLK90 = 1.33";
   attribute syn_tsu286: string;
   attribute syn_tsu286 of DEF_ARCH : architecture is " DATA_IN_1[70]->CLK = 1.335";
   attribute syn_tsu287: string;
   attribute syn_tsu287 of DEF_ARCH : architecture is " DATA_IN_1[70]->CLK90 = 1.33";
   attribute syn_tsu288: string;
   attribute syn_tsu288 of DEF_ARCH : architecture is " DATA_IN_1[71]->CLK = 1.335";
   attribute syn_tsu289: string;
   attribute syn_tsu289 of DEF_ARCH : architecture is " DATA_IN_1[71]->CLK90 = 1.33";
   attribute syn_tsu290: string;
   attribute syn_tsu290 of DEF_ARCH : architecture is " DATA_IN_1[72]->CLK = 1.335";
   attribute syn_tsu291: string;
   attribute syn_tsu291 of DEF_ARCH : architecture is " DATA_IN_1[72]->CLK90 = 1.33";
   attribute syn_tsu292: string;
   attribute syn_tsu292 of DEF_ARCH : architecture is " DATA_IN_1[73]->CLK = 1.335";
   attribute syn_tsu293: string;
   attribute syn_tsu293 of DEF_ARCH : architecture is " DATA_IN_1[73]->CLK90 = 1.33";
   attribute syn_tsu294: string;
   attribute syn_tsu294 of DEF_ARCH : architecture is " DATA_IN_1[74]->CLK = 1.335";
   attribute syn_tsu295: string;
   attribute syn_tsu295 of DEF_ARCH : architecture is " DATA_IN_1[74]->CLK90 = 1.33";
   attribute syn_tsu296: string;
   attribute syn_tsu296 of DEF_ARCH : architecture is " DATA_IN_1[75]->CLK = 1.335";
   attribute syn_tsu297: string;
   attribute syn_tsu297 of DEF_ARCH : architecture is " DATA_IN_1[75]->CLK90 = 1.33";
   attribute syn_tsu298: string;
   attribute syn_tsu298 of DEF_ARCH : architecture is " DATA_IN_1[76]->CLK = 1.335";
   attribute syn_tsu299: string;
   attribute syn_tsu299 of DEF_ARCH : architecture is " DATA_IN_1[76]->CLK90 = 1.33";
   attribute syn_tsu300: string;
   attribute syn_tsu300 of DEF_ARCH : architecture is " DATA_IN_1[77]->CLK = 1.335";
   attribute syn_tsu301: string;
   attribute syn_tsu301 of DEF_ARCH : architecture is " DATA_IN_1[77]->CLK90 = 1.33";
   attribute syn_tsu302: string;
   attribute syn_tsu302 of DEF_ARCH : architecture is " DATA_IN_1[78]->CLK = 1.335";
   attribute syn_tsu303: string;
   attribute syn_tsu303 of DEF_ARCH : architecture is " DATA_IN_1[78]->CLK90 = 1.33";
   attribute syn_tsu304: string;
   attribute syn_tsu304 of DEF_ARCH : architecture is " DATA_IN_1[79]->CLK = 1.335";
   attribute syn_tsu305: string;
   attribute syn_tsu305 of DEF_ARCH : architecture is " DATA_IN_1[79]->CLK90 = 1.33";
   attribute syn_tsu306: string;
   attribute syn_tsu306 of DEF_ARCH : architecture is " DATA_IN_1[7]->CLK = 1.335";
   attribute syn_tsu307: string;
   attribute syn_tsu307 of DEF_ARCH : architecture is " DATA_IN_1[7]->CLK90 = 1.33";
   attribute syn_tsu308: string;
   attribute syn_tsu308 of DEF_ARCH : architecture is " DATA_IN_1[80]->CLK = 1.335";
   attribute syn_tsu309: string;
   attribute syn_tsu309 of DEF_ARCH : architecture is " DATA_IN_1[80]->CLK90 = 1.33";
   attribute syn_tsu310: string;
   attribute syn_tsu310 of DEF_ARCH : architecture is " DATA_IN_1[81]->CLK = 1.335";
   attribute syn_tsu311: string;
   attribute syn_tsu311 of DEF_ARCH : architecture is " DATA_IN_1[81]->CLK90 = 1.33";
   attribute syn_tsu312: string;
   attribute syn_tsu312 of DEF_ARCH : architecture is " DATA_IN_1[82]->CLK = 1.335";
   attribute syn_tsu313: string;
   attribute syn_tsu313 of DEF_ARCH : architecture is " DATA_IN_1[82]->CLK90 = 1.33";
   attribute syn_tsu314: string;
   attribute syn_tsu314 of DEF_ARCH : architecture is " DATA_IN_1[83]->CLK = 1.335";
   attribute syn_tsu315: string;
   attribute syn_tsu315 of DEF_ARCH : architecture is " DATA_IN_1[83]->CLK90 = 1.33";
   attribute syn_tsu316: string;
   attribute syn_tsu316 of DEF_ARCH : architecture is " DATA_IN_1[84]->CLK = 1.335";
   attribute syn_tsu317: string;
   attribute syn_tsu317 of DEF_ARCH : architecture is " DATA_IN_1[84]->CLK90 = 1.33";
   attribute syn_tsu318: string;
   attribute syn_tsu318 of DEF_ARCH : architecture is " DATA_IN_1[85]->CLK = 1.335";
   attribute syn_tsu319: string;
   attribute syn_tsu319 of DEF_ARCH : architecture is " DATA_IN_1[85]->CLK90 = 1.33";
   attribute syn_tsu320: string;
   attribute syn_tsu320 of DEF_ARCH : architecture is " DATA_IN_1[86]->CLK = 1.335";
   attribute syn_tsu321: string;
   attribute syn_tsu321 of DEF_ARCH : architecture is " DATA_IN_1[86]->CLK90 = 1.33";
   attribute syn_tsu322: string;
   attribute syn_tsu322 of DEF_ARCH : architecture is " DATA_IN_1[87]->CLK = 1.335";
   attribute syn_tsu323: string;
   attribute syn_tsu323 of DEF_ARCH : architecture is " DATA_IN_1[87]->CLK90 = 1.33";
   attribute syn_tsu324: string;
   attribute syn_tsu324 of DEF_ARCH : architecture is " DATA_IN_1[88]->CLK = 1.335";
   attribute syn_tsu325: string;
   attribute syn_tsu325 of DEF_ARCH : architecture is " DATA_IN_1[88]->CLK90 = 1.33";
   attribute syn_tsu326: string;
   attribute syn_tsu326 of DEF_ARCH : architecture is " DATA_IN_1[89]->CLK = 1.335";
   attribute syn_tsu327: string;
   attribute syn_tsu327 of DEF_ARCH : architecture is " DATA_IN_1[89]->CLK90 = 1.33";
   attribute syn_tsu328: string;
   attribute syn_tsu328 of DEF_ARCH : architecture is " DATA_IN_1[8]->CLK = 1.335";
   attribute syn_tsu329: string;
   attribute syn_tsu329 of DEF_ARCH : architecture is " DATA_IN_1[8]->CLK90 = 1.33";
   attribute syn_tsu330: string;
   attribute syn_tsu330 of DEF_ARCH : architecture is " DATA_IN_1[90]->CLK = 1.335";
   attribute syn_tsu331: string;
   attribute syn_tsu331 of DEF_ARCH : architecture is " DATA_IN_1[90]->CLK90 = 1.33";
   attribute syn_tsu332: string;
   attribute syn_tsu332 of DEF_ARCH : architecture is " DATA_IN_1[91]->CLK = 1.335";
   attribute syn_tsu333: string;
   attribute syn_tsu333 of DEF_ARCH : architecture is " DATA_IN_1[91]->CLK90 = 1.33";
   attribute syn_tsu334: string;
   attribute syn_tsu334 of DEF_ARCH : architecture is " DATA_IN_1[92]->CLK = 1.335";
   attribute syn_tsu335: string;
   attribute syn_tsu335 of DEF_ARCH : architecture is " DATA_IN_1[92]->CLK90 = 1.33";
   attribute syn_tsu336: string;
   attribute syn_tsu336 of DEF_ARCH : architecture is " DATA_IN_1[93]->CLK = 1.335";
   attribute syn_tsu337: string;
   attribute syn_tsu337 of DEF_ARCH : architecture is " DATA_IN_1[93]->CLK90 = 1.33";
   attribute syn_tsu338: string;
   attribute syn_tsu338 of DEF_ARCH : architecture is " DATA_IN_1[94]->CLK = 1.335";
   attribute syn_tsu339: string;
   attribute syn_tsu339 of DEF_ARCH : architecture is " DATA_IN_1[94]->CLK90 = 1.33";
   attribute syn_tsu340: string;
   attribute syn_tsu340 of DEF_ARCH : architecture is " DATA_IN_1[95]->CLK = 1.335";
   attribute syn_tsu341: string;
   attribute syn_tsu341 of DEF_ARCH : architecture is " DATA_IN_1[95]->CLK90 = 1.33";
   attribute syn_tsu342: string;
   attribute syn_tsu342 of DEF_ARCH : architecture is " DATA_IN_1[96]->CLK = 1.335";
   attribute syn_tsu343: string;
   attribute syn_tsu343 of DEF_ARCH : architecture is " DATA_IN_1[96]->CLK90 = 1.33";
   attribute syn_tsu344: string;
   attribute syn_tsu344 of DEF_ARCH : architecture is " DATA_IN_1[97]->CLK = 1.335";
   attribute syn_tsu345: string;
   attribute syn_tsu345 of DEF_ARCH : architecture is " DATA_IN_1[97]->CLK90 = 1.33";
   attribute syn_tsu346: string;
   attribute syn_tsu346 of DEF_ARCH : architecture is " DATA_IN_1[98]->CLK = 1.335";
   attribute syn_tsu347: string;
   attribute syn_tsu347 of DEF_ARCH : architecture is " DATA_IN_1[98]->CLK90 = 1.33";
   attribute syn_tsu348: string;
   attribute syn_tsu348 of DEF_ARCH : architecture is " DATA_IN_1[99]->CLK = 1.335";
   attribute syn_tsu349: string;
   attribute syn_tsu349 of DEF_ARCH : architecture is " DATA_IN_1[99]->CLK90 = 1.33";
   attribute syn_tsu350: string;
   attribute syn_tsu350 of DEF_ARCH : architecture is " DATA_IN_1[9]->CLK = 1.335";
   attribute syn_tsu351: string;
   attribute syn_tsu351 of DEF_ARCH : architecture is " DATA_IN_1[9]->CLK90 = 1.33";
   attribute syn_tsu352: string;
   attribute syn_tsu352 of DEF_ARCH : architecture is " LATCH->CLK = 0.428";
   attribute syn_tsu353: string;
   attribute syn_tsu353 of DEF_ARCH : architecture is " LATCH->OUT_CLK = 0.428";
   attribute syn_tsu354: string;
   attribute syn_tsu354 of DEF_ARCH : architecture is " SEND_DATA_0->OUT_CLK = 1.147";
   attribute syn_tsu355: string;
   attribute syn_tsu355 of DEF_ARCH : architecture is " SEND_DATA_1->OUT_CLK = 1.148";
   attribute syn_tsu356: string;
   attribute syn_tsu356 of DEF_ARCH : architecture is " SHIFT_EN->BCO_CLK = 0.454";
   attribute syn_tsu357: string;
   attribute syn_tsu357 of DEF_ARCH : architecture is " SHIFT_IN->BCO_CLK = 0.428";
   attribute syn_tsu358: string;
   attribute syn_tsu358 of DEF_ARCH : architecture is " TEST_OUT[0]->CLK = 1.335";
   attribute syn_tsu359: string;
   attribute syn_tsu359 of DEF_ARCH : architecture is " TEST_OUT[0]->CLK90 = 1.33";
   attribute syn_tco0: string;
   attribute syn_tco0 of DEF_ARCH : architecture is " BCO_CLK->SHIFT_OUT = 0.550";
   attribute syn_tco1: string;
   attribute syn_tco1 of DEF_ARCH : architecture is " CLK->TEST_OUT[1] = 0.550";
   attribute syn_tco2: string;
   attribute syn_tco2 of DEF_ARCH : architecture is " CLK->TEST_OUT[2] = 0.550";
   attribute syn_tpd3: string;
   attribute syn_tpd3 of DEF_ARCH : architecture is " DATA_IN_1[103]->TEST_OUT[0] = 0.000";
   attribute syn_tco4: string;
   attribute syn_tco4 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_0[0] = 0.550";
   attribute syn_tco5: string;
   attribute syn_tco5 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_0[10] = 0.550";
   attribute syn_tco6: string;
   attribute syn_tco6 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_0[11] = 0.550";
   attribute syn_tco7: string;
   attribute syn_tco7 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_0[12] = 0.550";
   attribute syn_tco8: string;
   attribute syn_tco8 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_0[13] = 0.550";
   attribute syn_tco9: string;
   attribute syn_tco9 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_0[14] = 0.550";
   attribute syn_tco10: string;
   attribute syn_tco10 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_0[15] = 0.550";
   attribute syn_tco11: string;
   attribute syn_tco11 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_0[16] = 0.550";
   attribute syn_tco12: string;
   attribute syn_tco12 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_0[17] = 0.550";
   attribute syn_tco13: string;
   attribute syn_tco13 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_0[18] = 0.550";
   attribute syn_tco14: string;
   attribute syn_tco14 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_0[19] = 0.550";
   attribute syn_tco15: string;
   attribute syn_tco15 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_0[1] = 0.550";
   attribute syn_tco16: string;
   attribute syn_tco16 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_0[20] = 0.550";
   attribute syn_tco17: string;
   attribute syn_tco17 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_0[21] = 0.550";
   attribute syn_tco18: string;
   attribute syn_tco18 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_0[22] = 0.550";
   attribute syn_tco19: string;
   attribute syn_tco19 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_0[23] = 0.550";
   attribute syn_tco20: string;
   attribute syn_tco20 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_0[24] = 0.550";
   attribute syn_tco21: string;
   attribute syn_tco21 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_0[25] = 0.550";
   attribute syn_tco22: string;
   attribute syn_tco22 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_0[26] = 0.550";
   attribute syn_tco23: string;
   attribute syn_tco23 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_0[27] = 0.550";
   attribute syn_tco24: string;
   attribute syn_tco24 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_0[28] = 0.550";
   attribute syn_tco25: string;
   attribute syn_tco25 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_0[29] = 0.550";
   attribute syn_tco26: string;
   attribute syn_tco26 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_0[2] = 0.550";
   attribute syn_tco27: string;
   attribute syn_tco27 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_0[30] = 0.550";
   attribute syn_tco28: string;
   attribute syn_tco28 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_0[31] = 0.550";
   attribute syn_tco29: string;
   attribute syn_tco29 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_0[3] = 0.550";
   attribute syn_tco30: string;
   attribute syn_tco30 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_0[4] = 0.550";
   attribute syn_tco31: string;
   attribute syn_tco31 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_0[5] = 0.550";
   attribute syn_tco32: string;
   attribute syn_tco32 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_0[6] = 0.550";
   attribute syn_tco33: string;
   attribute syn_tco33 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_0[7] = 0.550";
   attribute syn_tco34: string;
   attribute syn_tco34 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_0[8] = 0.550";
   attribute syn_tco35: string;
   attribute syn_tco35 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_0[9] = 0.550";
   attribute syn_tco36: string;
   attribute syn_tco36 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_1[0] = 0.550";
   attribute syn_tco37: string;
   attribute syn_tco37 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_1[10] = 0.550";
   attribute syn_tco38: string;
   attribute syn_tco38 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_1[11] = 0.550";
   attribute syn_tco39: string;
   attribute syn_tco39 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_1[12] = 0.550";
   attribute syn_tco40: string;
   attribute syn_tco40 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_1[13] = 0.550";
   attribute syn_tco41: string;
   attribute syn_tco41 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_1[14] = 0.550";
   attribute syn_tco42: string;
   attribute syn_tco42 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_1[15] = 0.550";
   attribute syn_tco43: string;
   attribute syn_tco43 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_1[16] = 0.550";
   attribute syn_tco44: string;
   attribute syn_tco44 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_1[17] = 0.550";
   attribute syn_tco45: string;
   attribute syn_tco45 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_1[18] = 0.550";
   attribute syn_tco46: string;
   attribute syn_tco46 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_1[19] = 0.550";
   attribute syn_tco47: string;
   attribute syn_tco47 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_1[1] = 0.550";
   attribute syn_tco48: string;
   attribute syn_tco48 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_1[20] = 0.550";
   attribute syn_tco49: string;
   attribute syn_tco49 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_1[21] = 0.550";
   attribute syn_tco50: string;
   attribute syn_tco50 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_1[22] = 0.550";
   attribute syn_tco51: string;
   attribute syn_tco51 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_1[23] = 0.550";
   attribute syn_tco52: string;
   attribute syn_tco52 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_1[24] = 0.550";
   attribute syn_tco53: string;
   attribute syn_tco53 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_1[25] = 0.550";
   attribute syn_tco54: string;
   attribute syn_tco54 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_1[26] = 0.550";
   attribute syn_tco55: string;
   attribute syn_tco55 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_1[27] = 0.550";
   attribute syn_tco56: string;
   attribute syn_tco56 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_1[28] = 0.550";
   attribute syn_tco57: string;
   attribute syn_tco57 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_1[29] = 0.550";
   attribute syn_tco58: string;
   attribute syn_tco58 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_1[2] = 0.550";
   attribute syn_tco59: string;
   attribute syn_tco59 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_1[30] = 0.550";
   attribute syn_tco60: string;
   attribute syn_tco60 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_1[31] = 0.550";
   attribute syn_tco61: string;
   attribute syn_tco61 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_1[3] = 0.550";
   attribute syn_tco62: string;
   attribute syn_tco62 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_1[4] = 0.550";
   attribute syn_tco63: string;
   attribute syn_tco63 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_1[5] = 0.550";
   attribute syn_tco64: string;
   attribute syn_tco64 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_1[6] = 0.550";
   attribute syn_tco65: string;
   attribute syn_tco65 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_1[7] = 0.550";
   attribute syn_tco66: string;
   attribute syn_tco66 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_1[8] = 0.550";
   attribute syn_tco67: string;
   attribute syn_tco67 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_1[9] = 0.550";
   attribute syn_tco68: string;
   attribute syn_tco68 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_2[0] = 0.550";
   attribute syn_tco69: string;
   attribute syn_tco69 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_2[10] = 0.550";
   attribute syn_tco70: string;
   attribute syn_tco70 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_2[11] = 0.550";
   attribute syn_tco71: string;
   attribute syn_tco71 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_2[12] = 0.550";
   attribute syn_tco72: string;
   attribute syn_tco72 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_2[13] = 0.550";
   attribute syn_tco73: string;
   attribute syn_tco73 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_2[14] = 0.550";
   attribute syn_tco74: string;
   attribute syn_tco74 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_2[15] = 0.550";
   attribute syn_tco75: string;
   attribute syn_tco75 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_2[16] = 0.550";
   attribute syn_tco76: string;
   attribute syn_tco76 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_2[17] = 0.550";
   attribute syn_tco77: string;
   attribute syn_tco77 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_2[18] = 0.550";
   attribute syn_tco78: string;
   attribute syn_tco78 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_2[19] = 0.550";
   attribute syn_tco79: string;
   attribute syn_tco79 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_2[1] = 0.550";
   attribute syn_tco80: string;
   attribute syn_tco80 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_2[20] = 0.550";
   attribute syn_tco81: string;
   attribute syn_tco81 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_2[21] = 0.550";
   attribute syn_tco82: string;
   attribute syn_tco82 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_2[22] = 0.550";
   attribute syn_tco83: string;
   attribute syn_tco83 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_2[23] = 0.550";
   attribute syn_tco84: string;
   attribute syn_tco84 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_2[24] = 0.550";
   attribute syn_tco85: string;
   attribute syn_tco85 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_2[25] = 0.550";
   attribute syn_tco86: string;
   attribute syn_tco86 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_2[26] = 0.550";
   attribute syn_tco87: string;
   attribute syn_tco87 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_2[27] = 0.550";
   attribute syn_tco88: string;
   attribute syn_tco88 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_2[28] = 0.550";
   attribute syn_tco89: string;
   attribute syn_tco89 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_2[29] = 0.550";
   attribute syn_tco90: string;
   attribute syn_tco90 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_2[2] = 0.550";
   attribute syn_tco91: string;
   attribute syn_tco91 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_2[30] = 0.550";
   attribute syn_tco92: string;
   attribute syn_tco92 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_2[31] = 0.550";
   attribute syn_tco93: string;
   attribute syn_tco93 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_2[3] = 0.550";
   attribute syn_tco94: string;
   attribute syn_tco94 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_2[4] = 0.550";
   attribute syn_tco95: string;
   attribute syn_tco95 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_2[5] = 0.550";
   attribute syn_tco96: string;
   attribute syn_tco96 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_2[6] = 0.550";
   attribute syn_tco97: string;
   attribute syn_tco97 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_2[7] = 0.550";
   attribute syn_tco98: string;
   attribute syn_tco98 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_2[8] = 0.550";
   attribute syn_tco99: string;
   attribute syn_tco99 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_2[9] = 0.550";
   attribute syn_tco100: string;
   attribute syn_tco100 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_3[0] = 0.550";
   attribute syn_tco101: string;
   attribute syn_tco101 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_3[10] = 0.550";
   attribute syn_tco102: string;
   attribute syn_tco102 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_3[11] = 0.550";
   attribute syn_tco103: string;
   attribute syn_tco103 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_3[12] = 0.550";
   attribute syn_tco104: string;
   attribute syn_tco104 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_3[13] = 0.550";
   attribute syn_tco105: string;
   attribute syn_tco105 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_3[14] = 0.550";
   attribute syn_tco106: string;
   attribute syn_tco106 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_3[15] = 0.550";
   attribute syn_tco107: string;
   attribute syn_tco107 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_3[16] = 0.550";
   attribute syn_tco108: string;
   attribute syn_tco108 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_3[17] = 0.550";
   attribute syn_tco109: string;
   attribute syn_tco109 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_3[18] = 0.550";
   attribute syn_tco110: string;
   attribute syn_tco110 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_3[19] = 0.550";
   attribute syn_tco111: string;
   attribute syn_tco111 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_3[1] = 0.550";
   attribute syn_tco112: string;
   attribute syn_tco112 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_3[20] = 0.550";
   attribute syn_tco113: string;
   attribute syn_tco113 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_3[21] = 0.550";
   attribute syn_tco114: string;
   attribute syn_tco114 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_3[22] = 0.550";
   attribute syn_tco115: string;
   attribute syn_tco115 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_3[23] = 0.550";
   attribute syn_tco116: string;
   attribute syn_tco116 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_3[24] = 0.550";
   attribute syn_tco117: string;
   attribute syn_tco117 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_3[25] = 0.550";
   attribute syn_tco118: string;
   attribute syn_tco118 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_3[26] = 0.550";
   attribute syn_tco119: string;
   attribute syn_tco119 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_3[27] = 0.550";
   attribute syn_tco120: string;
   attribute syn_tco120 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_3[28] = 0.550";
   attribute syn_tco121: string;
   attribute syn_tco121 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_3[29] = 0.550";
   attribute syn_tco122: string;
   attribute syn_tco122 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_3[2] = 0.550";
   attribute syn_tco123: string;
   attribute syn_tco123 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_3[30] = 0.550";
   attribute syn_tco124: string;
   attribute syn_tco124 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_3[31] = 0.550";
   attribute syn_tco125: string;
   attribute syn_tco125 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_3[3] = 0.550";
   attribute syn_tco126: string;
   attribute syn_tco126 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_3[4] = 0.550";
   attribute syn_tco127: string;
   attribute syn_tco127 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_3[5] = 0.550";
   attribute syn_tco128: string;
   attribute syn_tco128 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_3[6] = 0.550";
   attribute syn_tco129: string;
   attribute syn_tco129 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_3[7] = 0.550";
   attribute syn_tco130: string;
   attribute syn_tco130 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_3[8] = 0.550";
   attribute syn_tco131: string;
   attribute syn_tco131 of DEF_ARCH : architecture is " OUT_CLK->DATA_OUT_3[9] = 0.550";
   attribute syn_tco132: string;
   attribute syn_tco132 of DEF_ARCH : architecture is " OUT_CLK->LSB[0] = 0.550";
   attribute syn_tco133: string;
   attribute syn_tco133 of DEF_ARCH : architecture is " OUT_CLK->LSB[1] = 0.550";
   attribute syn_tco134: string;
   attribute syn_tco134 of DEF_ARCH : architecture is " OUT_CLK->LSB[2] = 0.550";
   attribute syn_tco135: string;
   attribute syn_tco135 of DEF_ARCH : architecture is " OUT_CLK->LSB[3] = 0.550";
   attribute syn_tco136: string;
   attribute syn_tco136 of DEF_ARCH : architecture is " OUT_CLK->LSB[4] = 0.550";
   attribute syn_tco137: string;
   attribute syn_tco137 of DEF_ARCH : architecture is " OUT_CLK->LSB[5] = 0.550";
   attribute syn_tco138: string;
   attribute syn_tco138 of DEF_ARCH : architecture is " OUT_CLK->LSB[6] = 0.550";
   attribute syn_tco139: string;
   attribute syn_tco139 of DEF_ARCH : architecture is " OUT_CLK->LSB[7] = 0.550";
   attribute syn_tco140: string;
   attribute syn_tco140 of DEF_ARCH : architecture is " OUT_CLK->MSB[0] = 0.550";
   attribute syn_tco141: string;
   attribute syn_tco141 of DEF_ARCH : architecture is " OUT_CLK->MSB[1] = 0.550";
   attribute syn_tco142: string;
   attribute syn_tco142 of DEF_ARCH : architecture is " OUT_CLK->MSB[2] = 0.550";
   attribute syn_tco143: string;
   attribute syn_tco143 of DEF_ARCH : architecture is " OUT_CLK->MSB[3] = 0.550";
   attribute syn_tco144: string;
   attribute syn_tco144 of DEF_ARCH : architecture is " OUT_CLK->MSB[4] = 0.550";
   attribute syn_tco145: string;
   attribute syn_tco145 of DEF_ARCH : architecture is " OUT_CLK->MSB[5] = 0.550";
   attribute syn_tco146: string;
   attribute syn_tco146 of DEF_ARCH : architecture is " OUT_CLK->MSB[6] = 0.550";
   attribute syn_tco147: string;
   attribute syn_tco147 of DEF_ARCH : architecture is " OUT_CLK->MSB[7] = 0.550";
   attribute syn_tco148: string;
   attribute syn_tco148 of DEF_ARCH : architecture is " OUT_CLK->TEST_OUT[3] = 0.550";
   attribute syn_tco149: string;
   attribute syn_tco149 of DEF_ARCH : architecture is " OUT_CLK->TEST_OUT[4] = 0.550";
   attribute syn_tpd150: string;
   attribute syn_tpd150 of DEF_ARCH : architecture is " TEST_OUT[0]->DATA_IN_1[103] = 0.000";
   attribute black_box_pad_pin : string;
   attribute black_box_pad_pin of DEF_ARCH : architecture is "";

begin

end DEF_ARCH;
