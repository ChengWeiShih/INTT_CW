-- Version: 9.1 SP5 9.1.5.1

library ieee;
use ieee.std_logic_1164.all;
library proasic3e;
use proasic3e.all;

entity roc_block is

    port( RST         : in    std_logic;
          BCO_CLK     : in    std_logic;
          CLK         : in    std_logic;
          CLK90       : in    std_logic;
          OUT_CLK     : in    std_logic;
          LATCH       : in    std_logic;
          SEND_DATA_0 : in    std_logic;
          SEND_DATA_1 : in    std_logic;
          DATA_IN_0   : in    std_logic_vector(71 downto 0);
          DATA_IN_1   : in    std_logic_vector(103 downto 0);
          SHIFT_IN    : in    std_logic;
          SHIFT_EN    : in    std_logic;
          SHIFT_OUT   : out   std_logic;
          LSB         : out   std_logic_vector(7 downto 0);
          MSB         : out   std_logic_vector(7 downto 0);
          DATA_OUT_0  : out   std_logic_vector(31 downto 0);
          DATA_OUT_1  : out   std_logic_vector(31 downto 0);
          DATA_OUT_2  : out   std_logic_vector(31 downto 0);
          DATA_OUT_3  : out   std_logic_vector(31 downto 0);
          TEST_OUT    : out   std_logic_vector(7 downto 0)
        );

end roc_block;

architecture DEF_ARCH of roc_block is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component or_array
    port( CLK          : in    std_logic := 'U';
          RST          : in    std_logic := 'U';
          DATA_IN_0_0  : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_0_1  : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_0_2  : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_0_3  : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_0_4  : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_0_5  : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_0_6  : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_0_7  : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_0_8  : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_0_9  : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_0_26 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_0_27 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_0_28 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_0_29 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_0_30 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_0_31 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_0_32 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_0_33 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_0_34 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_0_35 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_0_36 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_0_37 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_0_38 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_0_39 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_0_40 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_0_41 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_0_42 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_0_43 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_0_44 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_0_45 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_0_46 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_0_47 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_0_48 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_0_49 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_0_50 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_0_51 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_0  : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_1  : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_2  : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_3  : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_4  : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_5  : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_6  : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_7  : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_8  : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_9  : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_10 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_11 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_12 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_13 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_14 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_15 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_16 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_17 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_18 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_19 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_20 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_21 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_22 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_23 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_24 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_25 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_26 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_27 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_28 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_29 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_30 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_31 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_32 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_33 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_34 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_35 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_36 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_37 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_38 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_39 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_40 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_41 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_42 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_43 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_44 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_45 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_46 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_47 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_48 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_49 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_50 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_IN_1_51 : in    std_logic_vector(25 downto 0) := (others => 'U');
          DATA_OUT_0_0 : out   std_logic_vector(25 downto 0);
          DATA_OUT_0_1 : out   std_logic_vector(25 downto 0);
          DATA_OUT_0_2 : out   std_logic_vector(25 downto 0);
          DATA_OUT_0_3 : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_0 : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_1 : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_2 : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_3 : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_4 : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_5 : out   std_logic_vector(25 downto 0)
        );
  end component;

  component decoder_array
    port( RST        : in    std_logic := 'U';
          CLK        : in    std_logic := 'U';
          CLR        : in    std_logic := 'U';
          DATA_OUT_0 : out   std_logic_vector(71 downto 0);
          DATA_OUT_1 : out   std_logic_vector(103 downto 0)
        );
  end component;

  component output_arbiter
    port( DATA_IN_0   : in    std_logic_vector(31 downto 0) := (others => 'U');
          DATA_IN_1   : in    std_logic_vector(31 downto 0) := (others => 'U');
          DATA_IN_2   : in    std_logic_vector(31 downto 0) := (others => 'U');
          DATA_IN_3   : in    std_logic_vector(31 downto 0) := (others => 'U');
          DATA_IN_4   : in    std_logic_vector(31 downto 0) := (others => 'U');
          DATA_IN_5   : in    std_logic_vector(31 downto 0) := (others => 'U');
          DATA_IN_6   : in    std_logic_vector(31 downto 0) := (others => 'U');
          DATA_IN_7   : in    std_logic_vector(31 downto 0) := (others => 'U');
          DATA_IN_8   : in    std_logic_vector(31 downto 0) := (others => 'U');
          DATA_IN_9   : in    std_logic_vector(31 downto 0) := (others => 'U');
          CLK         : in    std_logic := 'U';
          SEND_DATA_0 : in    std_logic := 'U';
          SEND_DATA_1 : in    std_logic := 'U';
          OUT_CLK     : in    std_logic := 'U';
          DATA_OUT_0  : out   std_logic_vector(31 downto 0);
          DATA_OUT_1  : out   std_logic_vector(31 downto 0);
          DATA_OUT_2  : out   std_logic_vector(31 downto 0);
          DATA_OUT_3  : out   std_logic_vector(31 downto 0);
          RST         : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component sync_block_logic
    port( RST        : in    std_logic := 'U';
          CLK        : in    std_logic := 'U';
          DATA_IN_0  : in    std_logic_vector(31 downto 0) := (others => 'U');
          DATA_IN_1  : in    std_logic_vector(31 downto 0) := (others => 'U');
          DATA_IN_2  : in    std_logic_vector(31 downto 0) := (others => 'U');
          DATA_IN_3  : in    std_logic_vector(31 downto 0) := (others => 'U');
          START      : in    std_logic := 'U';
          LSB        : out   std_logic_vector(7 downto 0);
          MSB        : out   std_logic_vector(7 downto 0);
          DATA_OUT_0 : out   std_logic_vector(31 downto 0);
          DATA_OUT_1 : out   std_logic_vector(31 downto 0);
          DATA_OUT_2 : out   std_logic_vector(31 downto 0);
          DATA_OUT_3 : out   std_logic_vector(31 downto 0)
        );
  end component;

  component pf_array
    port( RST        : in    std_logic := 'U';
          DATA_IN_0  : in    std_logic_vector(71 downto 0) := (others => 'U');
          DATA_IN_1  : in    std_logic_vector(103 downto 0) := (others => 'U');
          BCO_CLK    : in    std_logic := 'U';
          CLK        : in    std_logic := 'U';
          CLK90      : in    std_logic := 'U';
          LATCH      : in    std_logic := 'U';
          SHIFT_IN   : in    std_logic := 'U';
          SHIFT_EN   : in    std_logic := 'U';
          SHIFT_OUT  : out   std_logic;
          DATA_OUT_0 : out   std_logic_vector(71 downto 0);
          DATA_OUT_1 : out   std_logic_vector(103 downto 0)
        );
  end component;

  component deser_array
    port( RST           : in    std_logic := 'U';
          DATA_IN_0     : in    std_logic_vector(71 downto 0) := (others => 'U');
          DATA_IN_1     : in    std_logic_vector(103 downto 0) := (others => 'U');
          WRITE_EN_0    : in    std_logic_vector(71 downto 0) := (others => 'U');
          WRITE_EN_1    : in    std_logic_vector(103 downto 0) := (others => 'U');
          CLK           : in    std_logic := 'U';
          DATA_OUT_0_0  : out   std_logic_vector(25 downto 0);
          DATA_OUT_0_1  : out   std_logic_vector(25 downto 0);
          DATA_OUT_0_2  : out   std_logic_vector(25 downto 0);
          DATA_OUT_0_3  : out   std_logic_vector(25 downto 0);
          DATA_OUT_0_4  : out   std_logic_vector(25 downto 0);
          DATA_OUT_0_5  : out   std_logic_vector(25 downto 0);
          DATA_OUT_0_6  : out   std_logic_vector(25 downto 0);
          DATA_OUT_0_7  : out   std_logic_vector(25 downto 0);
          DATA_OUT_0_8  : out   std_logic_vector(25 downto 0);
          DATA_OUT_0_9  : out   std_logic_vector(25 downto 0);
          DATA_OUT_0_26 : out   std_logic_vector(25 downto 0);
          DATA_OUT_0_27 : out   std_logic_vector(25 downto 0);
          DATA_OUT_0_28 : out   std_logic_vector(25 downto 0);
          DATA_OUT_0_29 : out   std_logic_vector(25 downto 0);
          DATA_OUT_0_30 : out   std_logic_vector(25 downto 0);
          DATA_OUT_0_31 : out   std_logic_vector(25 downto 0);
          DATA_OUT_0_32 : out   std_logic_vector(25 downto 0);
          DATA_OUT_0_33 : out   std_logic_vector(25 downto 0);
          DATA_OUT_0_34 : out   std_logic_vector(25 downto 0);
          DATA_OUT_0_35 : out   std_logic_vector(25 downto 0);
          DATA_OUT_0_36 : out   std_logic_vector(25 downto 0);
          DATA_OUT_0_37 : out   std_logic_vector(25 downto 0);
          DATA_OUT_0_38 : out   std_logic_vector(25 downto 0);
          DATA_OUT_0_39 : out   std_logic_vector(25 downto 0);
          DATA_OUT_0_40 : out   std_logic_vector(25 downto 0);
          DATA_OUT_0_41 : out   std_logic_vector(25 downto 0);
          DATA_OUT_0_42 : out   std_logic_vector(25 downto 0);
          DATA_OUT_0_43 : out   std_logic_vector(25 downto 0);
          DATA_OUT_0_44 : out   std_logic_vector(25 downto 0);
          DATA_OUT_0_45 : out   std_logic_vector(25 downto 0);
          DATA_OUT_0_46 : out   std_logic_vector(25 downto 0);
          DATA_OUT_0_47 : out   std_logic_vector(25 downto 0);
          DATA_OUT_0_48 : out   std_logic_vector(25 downto 0);
          DATA_OUT_0_49 : out   std_logic_vector(25 downto 0);
          DATA_OUT_0_50 : out   std_logic_vector(25 downto 0);
          DATA_OUT_0_51 : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_0  : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_1  : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_2  : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_3  : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_4  : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_5  : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_6  : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_7  : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_8  : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_9  : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_10 : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_11 : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_12 : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_13 : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_14 : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_15 : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_16 : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_17 : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_18 : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_19 : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_20 : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_21 : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_22 : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_23 : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_24 : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_25 : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_26 : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_27 : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_28 : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_29 : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_30 : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_31 : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_32 : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_33 : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_34 : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_35 : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_36 : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_37 : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_38 : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_39 : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_40 : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_41 : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_42 : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_43 : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_44 : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_45 : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_46 : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_47 : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_48 : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_49 : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_50 : out   std_logic_vector(25 downto 0);
          DATA_OUT_1_51 : out   std_logic_vector(25 downto 0)
        );
  end component;

    signal \DATA_IN_1[103]\, \DATA_OUT_PF_1[103]\, 
        \DATA_OUT_1_51[0]\, \DATA_OUT_3_tmp[0]\, 
        \DATA_OUT_2_tmp[0]\, \GND\, \DATA_OUT_PF_0[0]\, 
        \DATA_OUT_PF_0[1]\, \DATA_OUT_PF_0[2]\, 
        \DATA_OUT_PF_0[3]\, \DATA_OUT_PF_0[4]\, 
        \DATA_OUT_PF_0[5]\, \DATA_OUT_PF_0[6]\, 
        \DATA_OUT_PF_0[7]\, \DATA_OUT_PF_0[8]\, 
        \DATA_OUT_PF_0[9]\, \DATA_OUT_PF_0[10]\, 
        \DATA_OUT_PF_0[11]\, \DATA_OUT_PF_0[12]\, 
        \DATA_OUT_PF_0[13]\, \DATA_OUT_PF_0[14]\, 
        \DATA_OUT_PF_0[15]\, \DATA_OUT_PF_0[16]\, 
        \DATA_OUT_PF_0[17]\, \DATA_OUT_PF_0[18]\, 
        \DATA_OUT_PF_0[19]\, \DATA_OUT_PF_0[20]\, 
        \DATA_OUT_PF_0[21]\, \DATA_OUT_PF_0[22]\, 
        \DATA_OUT_PF_0[23]\, \DATA_OUT_PF_0[24]\, 
        \DATA_OUT_PF_0[25]\, \DATA_OUT_PF_0[26]\, 
        \DATA_OUT_PF_0[27]\, \DATA_OUT_PF_0[28]\, 
        \DATA_OUT_PF_0[29]\, \DATA_OUT_PF_0[30]\, 
        \DATA_OUT_PF_0[31]\, \DATA_OUT_PF_0[32]\, 
        \DATA_OUT_PF_0[33]\, \DATA_OUT_PF_0[34]\, 
        \DATA_OUT_PF_0[35]\, \DATA_OUT_PF_0[36]\, 
        \DATA_OUT_PF_0[37]\, \DATA_OUT_PF_0[38]\, 
        \DATA_OUT_PF_0[39]\, \DATA_OUT_PF_0[40]\, 
        \DATA_OUT_PF_0[41]\, \DATA_OUT_PF_0[42]\, 
        \DATA_OUT_PF_0[43]\, \DATA_OUT_PF_0[44]\, 
        \DATA_OUT_PF_0[45]\, \DATA_OUT_PF_0[46]\, 
        \DATA_OUT_PF_0[47]\, \DATA_OUT_PF_0[48]\, 
        \DATA_OUT_PF_0[49]\, \DATA_OUT_PF_0[50]\, 
        \DATA_OUT_PF_0[51]\, \DATA_OUT_PF_0[52]\, 
        \DATA_OUT_PF_0[53]\, \DATA_OUT_PF_0[54]\, 
        \DATA_OUT_PF_0[55]\, \DATA_OUT_PF_0[56]\, 
        \DATA_OUT_PF_0[57]\, \DATA_OUT_PF_0[58]\, 
        \DATA_OUT_PF_0[59]\, \DATA_OUT_PF_0[60]\, 
        \DATA_OUT_PF_0[61]\, \DATA_OUT_PF_0[62]\, 
        \DATA_OUT_PF_0[63]\, \DATA_OUT_PF_0[64]\, 
        \DATA_OUT_PF_0[65]\, \DATA_OUT_PF_0[66]\, 
        \DATA_OUT_PF_0[67]\, \DATA_OUT_PF_0[68]\, 
        \DATA_OUT_PF_0[69]\, \DATA_OUT_PF_0[70]\, 
        \DATA_OUT_PF_0[71]\, \DATA_OUT_PF_1[0]\, 
        \DATA_OUT_PF_1[1]\, \DATA_OUT_PF_1[2]\, 
        \DATA_OUT_PF_1[3]\, \DATA_OUT_PF_1[4]\, 
        \DATA_OUT_PF_1[5]\, \DATA_OUT_PF_1[6]\, 
        \DATA_OUT_PF_1[7]\, \DATA_OUT_PF_1[8]\, 
        \DATA_OUT_PF_1[9]\, \DATA_OUT_PF_1[10]\, 
        \DATA_OUT_PF_1[11]\, \DATA_OUT_PF_1[12]\, 
        \DATA_OUT_PF_1[13]\, \DATA_OUT_PF_1[14]\, 
        \DATA_OUT_PF_1[15]\, \DATA_OUT_PF_1[16]\, 
        \DATA_OUT_PF_1[17]\, \DATA_OUT_PF_1[18]\, 
        \DATA_OUT_PF_1[19]\, \DATA_OUT_PF_1[20]\, 
        \DATA_OUT_PF_1[21]\, \DATA_OUT_PF_1[22]\, 
        \DATA_OUT_PF_1[23]\, \DATA_OUT_PF_1[24]\, 
        \DATA_OUT_PF_1[25]\, \DATA_OUT_PF_1[26]\, 
        \DATA_OUT_PF_1[27]\, \DATA_OUT_PF_1[28]\, 
        \DATA_OUT_PF_1[29]\, \DATA_OUT_PF_1[30]\, 
        \DATA_OUT_PF_1[31]\, \DATA_OUT_PF_1[32]\, 
        \DATA_OUT_PF_1[33]\, \DATA_OUT_PF_1[34]\, 
        \DATA_OUT_PF_1[35]\, \DATA_OUT_PF_1[36]\, 
        \DATA_OUT_PF_1[37]\, \DATA_OUT_PF_1[38]\, 
        \DATA_OUT_PF_1[39]\, \DATA_OUT_PF_1[40]\, 
        \DATA_OUT_PF_1[41]\, \DATA_OUT_PF_1[42]\, 
        \DATA_OUT_PF_1[43]\, \DATA_OUT_PF_1[44]\, 
        \DATA_OUT_PF_1[45]\, \DATA_OUT_PF_1[46]\, 
        \DATA_OUT_PF_1[47]\, \DATA_OUT_PF_1[48]\, 
        \DATA_OUT_PF_1[49]\, \DATA_OUT_PF_1[50]\, 
        \DATA_OUT_PF_1[51]\, \DATA_OUT_PF_1[52]\, 
        \DATA_OUT_PF_1[53]\, \DATA_OUT_PF_1[54]\, 
        \DATA_OUT_PF_1[55]\, \DATA_OUT_PF_1[56]\, 
        \DATA_OUT_PF_1[57]\, \DATA_OUT_PF_1[58]\, 
        \DATA_OUT_PF_1[59]\, \DATA_OUT_PF_1[60]\, 
        \DATA_OUT_PF_1[61]\, \DATA_OUT_PF_1[62]\, 
        \DATA_OUT_PF_1[63]\, \DATA_OUT_PF_1[64]\, 
        \DATA_OUT_PF_1[65]\, \DATA_OUT_PF_1[66]\, 
        \DATA_OUT_PF_1[67]\, \DATA_OUT_PF_1[68]\, 
        \DATA_OUT_PF_1[69]\, \DATA_OUT_PF_1[70]\, 
        \DATA_OUT_PF_1[71]\, \DATA_OUT_PF_1[72]\, 
        \DATA_OUT_PF_1[73]\, \DATA_OUT_PF_1[74]\, 
        \DATA_OUT_PF_1[75]\, \DATA_OUT_PF_1[76]\, 
        \DATA_OUT_PF_1[77]\, \DATA_OUT_PF_1[78]\, 
        \DATA_OUT_PF_1[79]\, \DATA_OUT_PF_1[80]\, 
        \DATA_OUT_PF_1[81]\, \DATA_OUT_PF_1[82]\, 
        \DATA_OUT_PF_1[83]\, \DATA_OUT_PF_1[84]\, 
        \DATA_OUT_PF_1[85]\, \DATA_OUT_PF_1[86]\, 
        \DATA_OUT_PF_1[87]\, \DATA_OUT_PF_1[88]\, 
        \DATA_OUT_PF_1[89]\, \DATA_OUT_PF_1[90]\, 
        \DATA_OUT_PF_1[91]\, \DATA_OUT_PF_1[92]\, 
        \DATA_OUT_PF_1[93]\, \DATA_OUT_PF_1[94]\, 
        \DATA_OUT_PF_1[95]\, \DATA_OUT_PF_1[96]\, 
        \DATA_OUT_PF_1[97]\, \DATA_OUT_PF_1[98]\, 
        \DATA_OUT_PF_1[99]\, \DATA_OUT_PF_1[100]\, 
        \DATA_OUT_PF_1[101]\, \DATA_OUT_PF_1[102]\, 
        \WRITE_EN_0[0]\, \WRITE_EN_0[1]\, \WRITE_EN_0[2]\, 
        \WRITE_EN_0[3]\, \WRITE_EN_0[4]\, \WRITE_EN_0[5]\, 
        \WRITE_EN_0[6]\, \WRITE_EN_0[7]\, \WRITE_EN_0[8]\, 
        \WRITE_EN_0[9]\, \WRITE_EN_0[10]\, \WRITE_EN_0[11]\, 
        \WRITE_EN_0[12]\, \WRITE_EN_0[13]\, \WRITE_EN_0[14]\, 
        \WRITE_EN_0[15]\, \WRITE_EN_0[16]\, \WRITE_EN_0[17]\, 
        \WRITE_EN_0[18]\, \WRITE_EN_0[19]\, \WRITE_EN_0[20]\, 
        \WRITE_EN_0[21]\, \WRITE_EN_0[22]\, \WRITE_EN_0[23]\, 
        \WRITE_EN_0[24]\, \WRITE_EN_0[25]\, \WRITE_EN_0[26]\, 
        \WRITE_EN_0[27]\, \WRITE_EN_0[28]\, \WRITE_EN_0[29]\, 
        \WRITE_EN_0[30]\, \WRITE_EN_0[31]\, \WRITE_EN_0[32]\, 
        \WRITE_EN_0[33]\, \WRITE_EN_0[34]\, \WRITE_EN_0[35]\, 
        \WRITE_EN_0[36]\, \WRITE_EN_0[37]\, \WRITE_EN_0[38]\, 
        \WRITE_EN_0[39]\, \WRITE_EN_0[40]\, \WRITE_EN_0[41]\, 
        \WRITE_EN_0[42]\, \WRITE_EN_0[43]\, \WRITE_EN_0[44]\, 
        \WRITE_EN_0[45]\, \WRITE_EN_0[46]\, \WRITE_EN_0[47]\, 
        \WRITE_EN_0[48]\, \WRITE_EN_0[49]\, \WRITE_EN_0[50]\, 
        \WRITE_EN_0[51]\, \WRITE_EN_0[52]\, \WRITE_EN_0[53]\, 
        \WRITE_EN_0[54]\, \WRITE_EN_0[55]\, \WRITE_EN_0[56]\, 
        \WRITE_EN_0[57]\, \WRITE_EN_0[58]\, \WRITE_EN_0[59]\, 
        \WRITE_EN_0[60]\, \WRITE_EN_0[61]\, \WRITE_EN_0[62]\, 
        \WRITE_EN_0[63]\, \WRITE_EN_0[64]\, \WRITE_EN_0[65]\, 
        \WRITE_EN_0[66]\, \WRITE_EN_0[67]\, \WRITE_EN_0[68]\, 
        \WRITE_EN_0[69]\, \WRITE_EN_0[70]\, \WRITE_EN_0[71]\, 
        \WRITE_EN_1[0]\, \WRITE_EN_1[1]\, \WRITE_EN_1[2]\, 
        \WRITE_EN_1[3]\, \WRITE_EN_1[4]\, \WRITE_EN_1[5]\, 
        \WRITE_EN_1[6]\, \WRITE_EN_1[7]\, \WRITE_EN_1[8]\, 
        \WRITE_EN_1[9]\, \WRITE_EN_1[10]\, \WRITE_EN_1[11]\, 
        \WRITE_EN_1[12]\, \WRITE_EN_1[13]\, \WRITE_EN_1[14]\, 
        \WRITE_EN_1[15]\, \WRITE_EN_1[16]\, \WRITE_EN_1[17]\, 
        \WRITE_EN_1[18]\, \WRITE_EN_1[19]\, \WRITE_EN_1[20]\, 
        \WRITE_EN_1[21]\, \WRITE_EN_1[22]\, \WRITE_EN_1[23]\, 
        \WRITE_EN_1[24]\, \WRITE_EN_1[25]\, \WRITE_EN_1[26]\, 
        \WRITE_EN_1[27]\, \WRITE_EN_1[28]\, \WRITE_EN_1[29]\, 
        \WRITE_EN_1[30]\, \WRITE_EN_1[31]\, \WRITE_EN_1[32]\, 
        \WRITE_EN_1[33]\, \WRITE_EN_1[34]\, \WRITE_EN_1[35]\, 
        \WRITE_EN_1[36]\, \WRITE_EN_1[37]\, \WRITE_EN_1[38]\, 
        \WRITE_EN_1[39]\, \WRITE_EN_1[40]\, \WRITE_EN_1[41]\, 
        \WRITE_EN_1[42]\, \WRITE_EN_1[43]\, \WRITE_EN_1[44]\, 
        \WRITE_EN_1[45]\, \WRITE_EN_1[46]\, \WRITE_EN_1[47]\, 
        \WRITE_EN_1[48]\, \WRITE_EN_1[49]\, \WRITE_EN_1[50]\, 
        \WRITE_EN_1[51]\, \WRITE_EN_1[52]\, \WRITE_EN_1[53]\, 
        \WRITE_EN_1[54]\, \WRITE_EN_1[55]\, \WRITE_EN_1[56]\, 
        \WRITE_EN_1[57]\, \WRITE_EN_1[58]\, \WRITE_EN_1[59]\, 
        \WRITE_EN_1[60]\, \WRITE_EN_1[61]\, \WRITE_EN_1[62]\, 
        \WRITE_EN_1[63]\, \WRITE_EN_1[64]\, \WRITE_EN_1[65]\, 
        \WRITE_EN_1[66]\, \WRITE_EN_1[67]\, \WRITE_EN_1[68]\, 
        \WRITE_EN_1[69]\, \WRITE_EN_1[70]\, \WRITE_EN_1[71]\, 
        \WRITE_EN_1[72]\, \WRITE_EN_1[73]\, \WRITE_EN_1[74]\, 
        \WRITE_EN_1[75]\, \WRITE_EN_1[76]\, \WRITE_EN_1[77]\, 
        \WRITE_EN_1[78]\, \WRITE_EN_1[79]\, \WRITE_EN_1[80]\, 
        \WRITE_EN_1[81]\, \WRITE_EN_1[82]\, \WRITE_EN_1[83]\, 
        \WRITE_EN_1[84]\, \WRITE_EN_1[85]\, \WRITE_EN_1[86]\, 
        \WRITE_EN_1[87]\, \WRITE_EN_1[88]\, \WRITE_EN_1[89]\, 
        \WRITE_EN_1[90]\, \WRITE_EN_1[91]\, \WRITE_EN_1[92]\, 
        \WRITE_EN_1[93]\, \WRITE_EN_1[94]\, \WRITE_EN_1[95]\, 
        \WRITE_EN_1[96]\, \WRITE_EN_1[97]\, \WRITE_EN_1[98]\, 
        \WRITE_EN_1[99]\, \WRITE_EN_1[100]\, \WRITE_EN_1[101]\, 
        \WRITE_EN_1[102]\, \WRITE_EN_1[103]\, \DATA_OUT_0_0[0]\, 
        \DATA_OUT_0_0[1]\, \DATA_OUT_0_0[2]\, \DATA_OUT_0_0[3]\, 
        \DATA_OUT_0_0[4]\, \DATA_OUT_0_0[5]\, \DATA_OUT_0_0[6]\, 
        \DATA_OUT_0_0[7]\, \DATA_OUT_0_0[8]\, \DATA_OUT_0_0[9]\, 
        \DATA_OUT_0_0[10]\, \DATA_OUT_0_0[11]\, 
        \DATA_OUT_0_0[12]\, \DATA_OUT_0_0[13]\, 
        \DATA_OUT_0_0[14]\, \DATA_OUT_0_0[15]\, 
        \DATA_OUT_0_0[16]\, \DATA_OUT_0_0[17]\, 
        \DATA_OUT_0_0[18]\, \DATA_OUT_0_0[19]\, 
        \DATA_OUT_0_0[20]\, \DATA_OUT_0_0[21]\, 
        \DATA_OUT_0_0[22]\, \DATA_OUT_0_0[23]\, 
        \DATA_OUT_0_0[24]\, \DATA_OUT_0_0[25]\, \DATA_OUT_0_1[0]\, 
        \DATA_OUT_0_1[1]\, \DATA_OUT_0_1[2]\, \DATA_OUT_0_1[3]\, 
        \DATA_OUT_0_1[4]\, \DATA_OUT_0_1[5]\, \DATA_OUT_0_1[6]\, 
        \DATA_OUT_0_1[7]\, \DATA_OUT_0_1[8]\, \DATA_OUT_0_1[9]\, 
        \DATA_OUT_0_1[10]\, \DATA_OUT_0_1[11]\, 
        \DATA_OUT_0_1[12]\, \DATA_OUT_0_1[13]\, 
        \DATA_OUT_0_1[14]\, \DATA_OUT_0_1[15]\, 
        \DATA_OUT_0_1[16]\, \DATA_OUT_0_1[17]\, 
        \DATA_OUT_0_1[18]\, \DATA_OUT_0_1[19]\, 
        \DATA_OUT_0_1[20]\, \DATA_OUT_0_1[21]\, 
        \DATA_OUT_0_1[22]\, \DATA_OUT_0_1[23]\, 
        \DATA_OUT_0_1[24]\, \DATA_OUT_0_1[25]\, \DATA_OUT_0_2[0]\, 
        \DATA_OUT_0_2[1]\, \DATA_OUT_0_2[2]\, \DATA_OUT_0_2[3]\, 
        \DATA_OUT_0_2[4]\, \DATA_OUT_0_2[5]\, \DATA_OUT_0_2[6]\, 
        \DATA_OUT_0_2[7]\, \DATA_OUT_0_2[8]\, \DATA_OUT_0_2[9]\, 
        \DATA_OUT_0_2[10]\, \DATA_OUT_0_2[11]\, 
        \DATA_OUT_0_2[12]\, \DATA_OUT_0_2[13]\, 
        \DATA_OUT_0_2[14]\, \DATA_OUT_0_2[15]\, 
        \DATA_OUT_0_2[16]\, \DATA_OUT_0_2[17]\, 
        \DATA_OUT_0_2[18]\, \DATA_OUT_0_2[19]\, 
        \DATA_OUT_0_2[20]\, \DATA_OUT_0_2[21]\, 
        \DATA_OUT_0_2[22]\, \DATA_OUT_0_2[23]\, 
        \DATA_OUT_0_2[24]\, \DATA_OUT_0_2[25]\, \DATA_OUT_0_3[0]\, 
        \DATA_OUT_0_3[1]\, \DATA_OUT_0_3[2]\, \DATA_OUT_0_3[3]\, 
        \DATA_OUT_0_3[4]\, \DATA_OUT_0_3[5]\, \DATA_OUT_0_3[6]\, 
        \DATA_OUT_0_3[7]\, \DATA_OUT_0_3[8]\, \DATA_OUT_0_3[9]\, 
        \DATA_OUT_0_3[10]\, \DATA_OUT_0_3[11]\, 
        \DATA_OUT_0_3[12]\, \DATA_OUT_0_3[13]\, 
        \DATA_OUT_0_3[14]\, \DATA_OUT_0_3[15]\, 
        \DATA_OUT_0_3[16]\, \DATA_OUT_0_3[17]\, 
        \DATA_OUT_0_3[18]\, \DATA_OUT_0_3[19]\, 
        \DATA_OUT_0_3[20]\, \DATA_OUT_0_3[21]\, 
        \DATA_OUT_0_3[22]\, \DATA_OUT_0_3[23]\, 
        \DATA_OUT_0_3[24]\, \DATA_OUT_0_3[25]\, \DATA_OUT_0_4[0]\, 
        \DATA_OUT_0_4[1]\, \DATA_OUT_0_4[2]\, \DATA_OUT_0_4[3]\, 
        \DATA_OUT_0_4[4]\, \DATA_OUT_0_4[5]\, \DATA_OUT_0_4[6]\, 
        \DATA_OUT_0_4[7]\, \DATA_OUT_0_4[8]\, \DATA_OUT_0_4[9]\, 
        \DATA_OUT_0_4[10]\, \DATA_OUT_0_4[11]\, 
        \DATA_OUT_0_4[12]\, \DATA_OUT_0_4[13]\, 
        \DATA_OUT_0_4[14]\, \DATA_OUT_0_4[15]\, 
        \DATA_OUT_0_4[16]\, \DATA_OUT_0_4[17]\, 
        \DATA_OUT_0_4[18]\, \DATA_OUT_0_4[19]\, 
        \DATA_OUT_0_4[20]\, \DATA_OUT_0_4[21]\, 
        \DATA_OUT_0_4[22]\, \DATA_OUT_0_4[23]\, 
        \DATA_OUT_0_4[24]\, \DATA_OUT_0_4[25]\, \DATA_OUT_0_5[0]\, 
        \DATA_OUT_0_5[1]\, \DATA_OUT_0_5[2]\, \DATA_OUT_0_5[3]\, 
        \DATA_OUT_0_5[4]\, \DATA_OUT_0_5[5]\, \DATA_OUT_0_5[6]\, 
        \DATA_OUT_0_5[7]\, \DATA_OUT_0_5[8]\, \DATA_OUT_0_5[9]\, 
        \DATA_OUT_0_5[10]\, \DATA_OUT_0_5[11]\, 
        \DATA_OUT_0_5[12]\, \DATA_OUT_0_5[13]\, 
        \DATA_OUT_0_5[14]\, \DATA_OUT_0_5[15]\, 
        \DATA_OUT_0_5[16]\, \DATA_OUT_0_5[17]\, 
        \DATA_OUT_0_5[18]\, \DATA_OUT_0_5[19]\, 
        \DATA_OUT_0_5[20]\, \DATA_OUT_0_5[21]\, 
        \DATA_OUT_0_5[22]\, \DATA_OUT_0_5[23]\, 
        \DATA_OUT_0_5[24]\, \DATA_OUT_0_5[25]\, \DATA_OUT_0_6[0]\, 
        \DATA_OUT_0_6[1]\, \DATA_OUT_0_6[2]\, \DATA_OUT_0_6[3]\, 
        \DATA_OUT_0_6[4]\, \DATA_OUT_0_6[5]\, \DATA_OUT_0_6[6]\, 
        \DATA_OUT_0_6[7]\, \DATA_OUT_0_6[8]\, \DATA_OUT_0_6[9]\, 
        \DATA_OUT_0_6[10]\, \DATA_OUT_0_6[11]\, 
        \DATA_OUT_0_6[12]\, \DATA_OUT_0_6[13]\, 
        \DATA_OUT_0_6[14]\, \DATA_OUT_0_6[15]\, 
        \DATA_OUT_0_6[16]\, \DATA_OUT_0_6[17]\, 
        \DATA_OUT_0_6[18]\, \DATA_OUT_0_6[19]\, 
        \DATA_OUT_0_6[20]\, \DATA_OUT_0_6[21]\, 
        \DATA_OUT_0_6[22]\, \DATA_OUT_0_6[23]\, 
        \DATA_OUT_0_6[24]\, \DATA_OUT_0_6[25]\, \DATA_OUT_0_7[0]\, 
        \DATA_OUT_0_7[1]\, \DATA_OUT_0_7[2]\, \DATA_OUT_0_7[3]\, 
        \DATA_OUT_0_7[4]\, \DATA_OUT_0_7[5]\, \DATA_OUT_0_7[6]\, 
        \DATA_OUT_0_7[7]\, \DATA_OUT_0_7[8]\, \DATA_OUT_0_7[9]\, 
        \DATA_OUT_0_7[10]\, \DATA_OUT_0_7[11]\, 
        \DATA_OUT_0_7[12]\, \DATA_OUT_0_7[13]\, 
        \DATA_OUT_0_7[14]\, \DATA_OUT_0_7[15]\, 
        \DATA_OUT_0_7[16]\, \DATA_OUT_0_7[17]\, 
        \DATA_OUT_0_7[18]\, \DATA_OUT_0_7[19]\, 
        \DATA_OUT_0_7[20]\, \DATA_OUT_0_7[21]\, 
        \DATA_OUT_0_7[22]\, \DATA_OUT_0_7[23]\, 
        \DATA_OUT_0_7[24]\, \DATA_OUT_0_7[25]\, \DATA_OUT_0_8[0]\, 
        \DATA_OUT_0_8[1]\, \DATA_OUT_0_8[2]\, \DATA_OUT_0_8[3]\, 
        \DATA_OUT_0_8[4]\, \DATA_OUT_0_8[5]\, \DATA_OUT_0_8[6]\, 
        \DATA_OUT_0_8[7]\, \DATA_OUT_0_8[8]\, \DATA_OUT_0_8[9]\, 
        \DATA_OUT_0_8[10]\, \DATA_OUT_0_8[11]\, 
        \DATA_OUT_0_8[12]\, \DATA_OUT_0_8[13]\, 
        \DATA_OUT_0_8[14]\, \DATA_OUT_0_8[15]\, 
        \DATA_OUT_0_8[16]\, \DATA_OUT_0_8[17]\, 
        \DATA_OUT_0_8[18]\, \DATA_OUT_0_8[19]\, 
        \DATA_OUT_0_8[20]\, \DATA_OUT_0_8[21]\, 
        \DATA_OUT_0_8[22]\, \DATA_OUT_0_8[23]\, 
        \DATA_OUT_0_8[24]\, \DATA_OUT_0_8[25]\, \DATA_OUT_0_9[0]\, 
        \DATA_OUT_0_9[1]\, \DATA_OUT_0_9[2]\, \DATA_OUT_0_9[3]\, 
        \DATA_OUT_0_9[4]\, \DATA_OUT_0_9[5]\, \DATA_OUT_0_9[6]\, 
        \DATA_OUT_0_9[7]\, \DATA_OUT_0_9[8]\, \DATA_OUT_0_9[9]\, 
        \DATA_OUT_0_9[10]\, \DATA_OUT_0_9[11]\, 
        \DATA_OUT_0_9[12]\, \DATA_OUT_0_9[13]\, 
        \DATA_OUT_0_9[14]\, \DATA_OUT_0_9[15]\, 
        \DATA_OUT_0_9[16]\, \DATA_OUT_0_9[17]\, 
        \DATA_OUT_0_9[18]\, \DATA_OUT_0_9[19]\, 
        \DATA_OUT_0_9[20]\, \DATA_OUT_0_9[21]\, 
        \DATA_OUT_0_9[22]\, \DATA_OUT_0_9[23]\, 
        \DATA_OUT_0_9[24]\, \DATA_OUT_0_9[25]\, 
        \DATA_OUT_0_26[0]\, \DATA_OUT_0_26[1]\, 
        \DATA_OUT_0_26[2]\, \DATA_OUT_0_26[3]\, 
        \DATA_OUT_0_26[4]\, \DATA_OUT_0_26[5]\, 
        \DATA_OUT_0_26[6]\, \DATA_OUT_0_26[7]\, 
        \DATA_OUT_0_26[8]\, \DATA_OUT_0_26[9]\, 
        \DATA_OUT_0_26[10]\, \DATA_OUT_0_26[11]\, 
        \DATA_OUT_0_26[12]\, \DATA_OUT_0_26[13]\, 
        \DATA_OUT_0_26[14]\, \DATA_OUT_0_26[15]\, 
        \DATA_OUT_0_26[16]\, \DATA_OUT_0_26[17]\, 
        \DATA_OUT_0_26[18]\, \DATA_OUT_0_26[19]\, 
        \DATA_OUT_0_26[20]\, \DATA_OUT_0_26[21]\, 
        \DATA_OUT_0_26[22]\, \DATA_OUT_0_26[23]\, 
        \DATA_OUT_0_26[24]\, \DATA_OUT_0_26[25]\, 
        \DATA_OUT_0_27[0]\, \DATA_OUT_0_27[1]\, 
        \DATA_OUT_0_27[2]\, \DATA_OUT_0_27[3]\, 
        \DATA_OUT_0_27[4]\, \DATA_OUT_0_27[5]\, 
        \DATA_OUT_0_27[6]\, \DATA_OUT_0_27[7]\, 
        \DATA_OUT_0_27[8]\, \DATA_OUT_0_27[9]\, 
        \DATA_OUT_0_27[10]\, \DATA_OUT_0_27[11]\, 
        \DATA_OUT_0_27[12]\, \DATA_OUT_0_27[13]\, 
        \DATA_OUT_0_27[14]\, \DATA_OUT_0_27[15]\, 
        \DATA_OUT_0_27[16]\, \DATA_OUT_0_27[17]\, 
        \DATA_OUT_0_27[18]\, \DATA_OUT_0_27[19]\, 
        \DATA_OUT_0_27[20]\, \DATA_OUT_0_27[21]\, 
        \DATA_OUT_0_27[22]\, \DATA_OUT_0_27[23]\, 
        \DATA_OUT_0_27[24]\, \DATA_OUT_0_27[25]\, 
        \DATA_OUT_0_28[0]\, \DATA_OUT_0_28[1]\, 
        \DATA_OUT_0_28[2]\, \DATA_OUT_0_28[3]\, 
        \DATA_OUT_0_28[4]\, \DATA_OUT_0_28[5]\, 
        \DATA_OUT_0_28[6]\, \DATA_OUT_0_28[7]\, 
        \DATA_OUT_0_28[8]\, \DATA_OUT_0_28[9]\, 
        \DATA_OUT_0_28[10]\, \DATA_OUT_0_28[11]\, 
        \DATA_OUT_0_28[12]\, \DATA_OUT_0_28[13]\, 
        \DATA_OUT_0_28[14]\, \DATA_OUT_0_28[15]\, 
        \DATA_OUT_0_28[16]\, \DATA_OUT_0_28[17]\, 
        \DATA_OUT_0_28[18]\, \DATA_OUT_0_28[19]\, 
        \DATA_OUT_0_28[20]\, \DATA_OUT_0_28[21]\, 
        \DATA_OUT_0_28[22]\, \DATA_OUT_0_28[23]\, 
        \DATA_OUT_0_28[24]\, \DATA_OUT_0_28[25]\, 
        \DATA_OUT_0_29[0]\, \DATA_OUT_0_29[1]\, 
        \DATA_OUT_0_29[2]\, \DATA_OUT_0_29[3]\, 
        \DATA_OUT_0_29[4]\, \DATA_OUT_0_29[5]\, 
        \DATA_OUT_0_29[6]\, \DATA_OUT_0_29[7]\, 
        \DATA_OUT_0_29[8]\, \DATA_OUT_0_29[9]\, 
        \DATA_OUT_0_29[10]\, \DATA_OUT_0_29[11]\, 
        \DATA_OUT_0_29[12]\, \DATA_OUT_0_29[13]\, 
        \DATA_OUT_0_29[14]\, \DATA_OUT_0_29[15]\, 
        \DATA_OUT_0_29[16]\, \DATA_OUT_0_29[17]\, 
        \DATA_OUT_0_29[18]\, \DATA_OUT_0_29[19]\, 
        \DATA_OUT_0_29[20]\, \DATA_OUT_0_29[21]\, 
        \DATA_OUT_0_29[22]\, \DATA_OUT_0_29[23]\, 
        \DATA_OUT_0_29[24]\, \DATA_OUT_0_29[25]\, 
        \DATA_OUT_0_30[0]\, \DATA_OUT_0_30[1]\, 
        \DATA_OUT_0_30[2]\, \DATA_OUT_0_30[3]\, 
        \DATA_OUT_0_30[4]\, \DATA_OUT_0_30[5]\, 
        \DATA_OUT_0_30[6]\, \DATA_OUT_0_30[7]\, 
        \DATA_OUT_0_30[8]\, \DATA_OUT_0_30[9]\, 
        \DATA_OUT_0_30[10]\, \DATA_OUT_0_30[11]\, 
        \DATA_OUT_0_30[12]\, \DATA_OUT_0_30[13]\, 
        \DATA_OUT_0_30[14]\, \DATA_OUT_0_30[15]\, 
        \DATA_OUT_0_30[16]\, \DATA_OUT_0_30[17]\, 
        \DATA_OUT_0_30[18]\, \DATA_OUT_0_30[19]\, 
        \DATA_OUT_0_30[20]\, \DATA_OUT_0_30[21]\, 
        \DATA_OUT_0_30[22]\, \DATA_OUT_0_30[23]\, 
        \DATA_OUT_0_30[24]\, \DATA_OUT_0_30[25]\, 
        \DATA_OUT_0_31[0]\, \DATA_OUT_0_31[1]\, 
        \DATA_OUT_0_31[2]\, \DATA_OUT_0_31[3]\, 
        \DATA_OUT_0_31[4]\, \DATA_OUT_0_31[5]\, 
        \DATA_OUT_0_31[6]\, \DATA_OUT_0_31[7]\, 
        \DATA_OUT_0_31[8]\, \DATA_OUT_0_31[9]\, 
        \DATA_OUT_0_31[10]\, \DATA_OUT_0_31[11]\, 
        \DATA_OUT_0_31[12]\, \DATA_OUT_0_31[13]\, 
        \DATA_OUT_0_31[14]\, \DATA_OUT_0_31[15]\, 
        \DATA_OUT_0_31[16]\, \DATA_OUT_0_31[17]\, 
        \DATA_OUT_0_31[18]\, \DATA_OUT_0_31[19]\, 
        \DATA_OUT_0_31[20]\, \DATA_OUT_0_31[21]\, 
        \DATA_OUT_0_31[22]\, \DATA_OUT_0_31[23]\, 
        \DATA_OUT_0_31[24]\, \DATA_OUT_0_31[25]\, 
        \DATA_OUT_0_32[0]\, \DATA_OUT_0_32[1]\, 
        \DATA_OUT_0_32[2]\, \DATA_OUT_0_32[3]\, 
        \DATA_OUT_0_32[4]\, \DATA_OUT_0_32[5]\, 
        \DATA_OUT_0_32[6]\, \DATA_OUT_0_32[7]\, 
        \DATA_OUT_0_32[8]\, \DATA_OUT_0_32[9]\, 
        \DATA_OUT_0_32[10]\, \DATA_OUT_0_32[11]\, 
        \DATA_OUT_0_32[12]\, \DATA_OUT_0_32[13]\, 
        \DATA_OUT_0_32[14]\, \DATA_OUT_0_32[15]\, 
        \DATA_OUT_0_32[16]\, \DATA_OUT_0_32[17]\, 
        \DATA_OUT_0_32[18]\, \DATA_OUT_0_32[19]\, 
        \DATA_OUT_0_32[20]\, \DATA_OUT_0_32[21]\, 
        \DATA_OUT_0_32[22]\, \DATA_OUT_0_32[23]\, 
        \DATA_OUT_0_32[24]\, \DATA_OUT_0_32[25]\, 
        \DATA_OUT_0_33[0]\, \DATA_OUT_0_33[1]\, 
        \DATA_OUT_0_33[2]\, \DATA_OUT_0_33[3]\, 
        \DATA_OUT_0_33[4]\, \DATA_OUT_0_33[5]\, 
        \DATA_OUT_0_33[6]\, \DATA_OUT_0_33[7]\, 
        \DATA_OUT_0_33[8]\, \DATA_OUT_0_33[9]\, 
        \DATA_OUT_0_33[10]\, \DATA_OUT_0_33[11]\, 
        \DATA_OUT_0_33[12]\, \DATA_OUT_0_33[13]\, 
        \DATA_OUT_0_33[14]\, \DATA_OUT_0_33[15]\, 
        \DATA_OUT_0_33[16]\, \DATA_OUT_0_33[17]\, 
        \DATA_OUT_0_33[18]\, \DATA_OUT_0_33[19]\, 
        \DATA_OUT_0_33[20]\, \DATA_OUT_0_33[21]\, 
        \DATA_OUT_0_33[22]\, \DATA_OUT_0_33[23]\, 
        \DATA_OUT_0_33[24]\, \DATA_OUT_0_33[25]\, 
        \DATA_OUT_0_34[0]\, \DATA_OUT_0_34[1]\, 
        \DATA_OUT_0_34[2]\, \DATA_OUT_0_34[3]\, 
        \DATA_OUT_0_34[4]\, \DATA_OUT_0_34[5]\, 
        \DATA_OUT_0_34[6]\, \DATA_OUT_0_34[7]\, 
        \DATA_OUT_0_34[8]\, \DATA_OUT_0_34[9]\, 
        \DATA_OUT_0_34[10]\, \DATA_OUT_0_34[11]\, 
        \DATA_OUT_0_34[12]\, \DATA_OUT_0_34[13]\, 
        \DATA_OUT_0_34[14]\, \DATA_OUT_0_34[15]\, 
        \DATA_OUT_0_34[16]\, \DATA_OUT_0_34[17]\, 
        \DATA_OUT_0_34[18]\, \DATA_OUT_0_34[19]\, 
        \DATA_OUT_0_34[20]\, \DATA_OUT_0_34[21]\, 
        \DATA_OUT_0_34[22]\, \DATA_OUT_0_34[23]\, 
        \DATA_OUT_0_34[24]\, \DATA_OUT_0_34[25]\, 
        \DATA_OUT_0_35[0]\, \DATA_OUT_0_35[1]\, 
        \DATA_OUT_0_35[2]\, \DATA_OUT_0_35[3]\, 
        \DATA_OUT_0_35[4]\, \DATA_OUT_0_35[5]\, 
        \DATA_OUT_0_35[6]\, \DATA_OUT_0_35[7]\, 
        \DATA_OUT_0_35[8]\, \DATA_OUT_0_35[9]\, 
        \DATA_OUT_0_35[10]\, \DATA_OUT_0_35[11]\, 
        \DATA_OUT_0_35[12]\, \DATA_OUT_0_35[13]\, 
        \DATA_OUT_0_35[14]\, \DATA_OUT_0_35[15]\, 
        \DATA_OUT_0_35[16]\, \DATA_OUT_0_35[17]\, 
        \DATA_OUT_0_35[18]\, \DATA_OUT_0_35[19]\, 
        \DATA_OUT_0_35[20]\, \DATA_OUT_0_35[21]\, 
        \DATA_OUT_0_35[22]\, \DATA_OUT_0_35[23]\, 
        \DATA_OUT_0_35[24]\, \DATA_OUT_0_35[25]\, 
        \DATA_OUT_0_36[0]\, \DATA_OUT_0_36[1]\, 
        \DATA_OUT_0_36[2]\, \DATA_OUT_0_36[3]\, 
        \DATA_OUT_0_36[4]\, \DATA_OUT_0_36[5]\, 
        \DATA_OUT_0_36[6]\, \DATA_OUT_0_36[7]\, 
        \DATA_OUT_0_36[8]\, \DATA_OUT_0_36[9]\, 
        \DATA_OUT_0_36[10]\, \DATA_OUT_0_36[11]\, 
        \DATA_OUT_0_36[12]\, \DATA_OUT_0_36[13]\, 
        \DATA_OUT_0_36[14]\, \DATA_OUT_0_36[15]\, 
        \DATA_OUT_0_36[16]\, \DATA_OUT_0_36[17]\, 
        \DATA_OUT_0_36[18]\, \DATA_OUT_0_36[19]\, 
        \DATA_OUT_0_36[20]\, \DATA_OUT_0_36[21]\, 
        \DATA_OUT_0_36[22]\, \DATA_OUT_0_36[23]\, 
        \DATA_OUT_0_36[24]\, \DATA_OUT_0_36[25]\, 
        \DATA_OUT_0_37[0]\, \DATA_OUT_0_37[1]\, 
        \DATA_OUT_0_37[2]\, \DATA_OUT_0_37[3]\, 
        \DATA_OUT_0_37[4]\, \DATA_OUT_0_37[5]\, 
        \DATA_OUT_0_37[6]\, \DATA_OUT_0_37[7]\, 
        \DATA_OUT_0_37[8]\, \DATA_OUT_0_37[9]\, 
        \DATA_OUT_0_37[10]\, \DATA_OUT_0_37[11]\, 
        \DATA_OUT_0_37[12]\, \DATA_OUT_0_37[13]\, 
        \DATA_OUT_0_37[14]\, \DATA_OUT_0_37[15]\, 
        \DATA_OUT_0_37[16]\, \DATA_OUT_0_37[17]\, 
        \DATA_OUT_0_37[18]\, \DATA_OUT_0_37[19]\, 
        \DATA_OUT_0_37[20]\, \DATA_OUT_0_37[21]\, 
        \DATA_OUT_0_37[22]\, \DATA_OUT_0_37[23]\, 
        \DATA_OUT_0_37[24]\, \DATA_OUT_0_37[25]\, 
        \DATA_OUT_0_38[0]\, \DATA_OUT_0_38[1]\, 
        \DATA_OUT_0_38[2]\, \DATA_OUT_0_38[3]\, 
        \DATA_OUT_0_38[4]\, \DATA_OUT_0_38[5]\, 
        \DATA_OUT_0_38[6]\, \DATA_OUT_0_38[7]\, 
        \DATA_OUT_0_38[8]\, \DATA_OUT_0_38[9]\, 
        \DATA_OUT_0_38[10]\, \DATA_OUT_0_38[11]\, 
        \DATA_OUT_0_38[12]\, \DATA_OUT_0_38[13]\, 
        \DATA_OUT_0_38[14]\, \DATA_OUT_0_38[15]\, 
        \DATA_OUT_0_38[16]\, \DATA_OUT_0_38[17]\, 
        \DATA_OUT_0_38[18]\, \DATA_OUT_0_38[19]\, 
        \DATA_OUT_0_38[20]\, \DATA_OUT_0_38[21]\, 
        \DATA_OUT_0_38[22]\, \DATA_OUT_0_38[23]\, 
        \DATA_OUT_0_38[24]\, \DATA_OUT_0_38[25]\, 
        \DATA_OUT_0_39[0]\, \DATA_OUT_0_39[1]\, 
        \DATA_OUT_0_39[2]\, \DATA_OUT_0_39[3]\, 
        \DATA_OUT_0_39[4]\, \DATA_OUT_0_39[5]\, 
        \DATA_OUT_0_39[6]\, \DATA_OUT_0_39[7]\, 
        \DATA_OUT_0_39[8]\, \DATA_OUT_0_39[9]\, 
        \DATA_OUT_0_39[10]\, \DATA_OUT_0_39[11]\, 
        \DATA_OUT_0_39[12]\, \DATA_OUT_0_39[13]\, 
        \DATA_OUT_0_39[14]\, \DATA_OUT_0_39[15]\, 
        \DATA_OUT_0_39[16]\, \DATA_OUT_0_39[17]\, 
        \DATA_OUT_0_39[18]\, \DATA_OUT_0_39[19]\, 
        \DATA_OUT_0_39[20]\, \DATA_OUT_0_39[21]\, 
        \DATA_OUT_0_39[22]\, \DATA_OUT_0_39[23]\, 
        \DATA_OUT_0_39[24]\, \DATA_OUT_0_39[25]\, 
        \DATA_OUT_0_40[0]\, \DATA_OUT_0_40[1]\, 
        \DATA_OUT_0_40[2]\, \DATA_OUT_0_40[3]\, 
        \DATA_OUT_0_40[4]\, \DATA_OUT_0_40[5]\, 
        \DATA_OUT_0_40[6]\, \DATA_OUT_0_40[7]\, 
        \DATA_OUT_0_40[8]\, \DATA_OUT_0_40[9]\, 
        \DATA_OUT_0_40[10]\, \DATA_OUT_0_40[11]\, 
        \DATA_OUT_0_40[12]\, \DATA_OUT_0_40[13]\, 
        \DATA_OUT_0_40[14]\, \DATA_OUT_0_40[15]\, 
        \DATA_OUT_0_40[16]\, \DATA_OUT_0_40[17]\, 
        \DATA_OUT_0_40[18]\, \DATA_OUT_0_40[19]\, 
        \DATA_OUT_0_40[20]\, \DATA_OUT_0_40[21]\, 
        \DATA_OUT_0_40[22]\, \DATA_OUT_0_40[23]\, 
        \DATA_OUT_0_40[24]\, \DATA_OUT_0_40[25]\, 
        \DATA_OUT_0_41[0]\, \DATA_OUT_0_41[1]\, 
        \DATA_OUT_0_41[2]\, \DATA_OUT_0_41[3]\, 
        \DATA_OUT_0_41[4]\, \DATA_OUT_0_41[5]\, 
        \DATA_OUT_0_41[6]\, \DATA_OUT_0_41[7]\, 
        \DATA_OUT_0_41[8]\, \DATA_OUT_0_41[9]\, 
        \DATA_OUT_0_41[10]\, \DATA_OUT_0_41[11]\, 
        \DATA_OUT_0_41[12]\, \DATA_OUT_0_41[13]\, 
        \DATA_OUT_0_41[14]\, \DATA_OUT_0_41[15]\, 
        \DATA_OUT_0_41[16]\, \DATA_OUT_0_41[17]\, 
        \DATA_OUT_0_41[18]\, \DATA_OUT_0_41[19]\, 
        \DATA_OUT_0_41[20]\, \DATA_OUT_0_41[21]\, 
        \DATA_OUT_0_41[22]\, \DATA_OUT_0_41[23]\, 
        \DATA_OUT_0_41[24]\, \DATA_OUT_0_41[25]\, 
        \DATA_OUT_0_42[0]\, \DATA_OUT_0_42[1]\, 
        \DATA_OUT_0_42[2]\, \DATA_OUT_0_42[3]\, 
        \DATA_OUT_0_42[4]\, \DATA_OUT_0_42[5]\, 
        \DATA_OUT_0_42[6]\, \DATA_OUT_0_42[7]\, 
        \DATA_OUT_0_42[8]\, \DATA_OUT_0_42[9]\, 
        \DATA_OUT_0_42[10]\, \DATA_OUT_0_42[11]\, 
        \DATA_OUT_0_42[12]\, \DATA_OUT_0_42[13]\, 
        \DATA_OUT_0_42[14]\, \DATA_OUT_0_42[15]\, 
        \DATA_OUT_0_42[16]\, \DATA_OUT_0_42[17]\, 
        \DATA_OUT_0_42[18]\, \DATA_OUT_0_42[19]\, 
        \DATA_OUT_0_42[20]\, \DATA_OUT_0_42[21]\, 
        \DATA_OUT_0_42[22]\, \DATA_OUT_0_42[23]\, 
        \DATA_OUT_0_42[24]\, \DATA_OUT_0_42[25]\, 
        \DATA_OUT_0_43[0]\, \DATA_OUT_0_43[1]\, 
        \DATA_OUT_0_43[2]\, \DATA_OUT_0_43[3]\, 
        \DATA_OUT_0_43[4]\, \DATA_OUT_0_43[5]\, 
        \DATA_OUT_0_43[6]\, \DATA_OUT_0_43[7]\, 
        \DATA_OUT_0_43[8]\, \DATA_OUT_0_43[9]\, 
        \DATA_OUT_0_43[10]\, \DATA_OUT_0_43[11]\, 
        \DATA_OUT_0_43[12]\, \DATA_OUT_0_43[13]\, 
        \DATA_OUT_0_43[14]\, \DATA_OUT_0_43[15]\, 
        \DATA_OUT_0_43[16]\, \DATA_OUT_0_43[17]\, 
        \DATA_OUT_0_43[18]\, \DATA_OUT_0_43[19]\, 
        \DATA_OUT_0_43[20]\, \DATA_OUT_0_43[21]\, 
        \DATA_OUT_0_43[22]\, \DATA_OUT_0_43[23]\, 
        \DATA_OUT_0_43[24]\, \DATA_OUT_0_43[25]\, 
        \DATA_OUT_0_44[0]\, \DATA_OUT_0_44[1]\, 
        \DATA_OUT_0_44[2]\, \DATA_OUT_0_44[3]\, 
        \DATA_OUT_0_44[4]\, \DATA_OUT_0_44[5]\, 
        \DATA_OUT_0_44[6]\, \DATA_OUT_0_44[7]\, 
        \DATA_OUT_0_44[8]\, \DATA_OUT_0_44[9]\, 
        \DATA_OUT_0_44[10]\, \DATA_OUT_0_44[11]\, 
        \DATA_OUT_0_44[12]\, \DATA_OUT_0_44[13]\, 
        \DATA_OUT_0_44[14]\, \DATA_OUT_0_44[15]\, 
        \DATA_OUT_0_44[16]\, \DATA_OUT_0_44[17]\, 
        \DATA_OUT_0_44[18]\, \DATA_OUT_0_44[19]\, 
        \DATA_OUT_0_44[20]\, \DATA_OUT_0_44[21]\, 
        \DATA_OUT_0_44[22]\, \DATA_OUT_0_44[23]\, 
        \DATA_OUT_0_44[24]\, \DATA_OUT_0_44[25]\, 
        \DATA_OUT_0_45[0]\, \DATA_OUT_0_45[1]\, 
        \DATA_OUT_0_45[2]\, \DATA_OUT_0_45[3]\, 
        \DATA_OUT_0_45[4]\, \DATA_OUT_0_45[5]\, 
        \DATA_OUT_0_45[6]\, \DATA_OUT_0_45[7]\, 
        \DATA_OUT_0_45[8]\, \DATA_OUT_0_45[9]\, 
        \DATA_OUT_0_45[10]\, \DATA_OUT_0_45[11]\, 
        \DATA_OUT_0_45[12]\, \DATA_OUT_0_45[13]\, 
        \DATA_OUT_0_45[14]\, \DATA_OUT_0_45[15]\, 
        \DATA_OUT_0_45[16]\, \DATA_OUT_0_45[17]\, 
        \DATA_OUT_0_45[18]\, \DATA_OUT_0_45[19]\, 
        \DATA_OUT_0_45[20]\, \DATA_OUT_0_45[21]\, 
        \DATA_OUT_0_45[22]\, \DATA_OUT_0_45[23]\, 
        \DATA_OUT_0_45[24]\, \DATA_OUT_0_45[25]\, 
        \DATA_OUT_0_46[0]\, \DATA_OUT_0_46[1]\, 
        \DATA_OUT_0_46[2]\, \DATA_OUT_0_46[3]\, 
        \DATA_OUT_0_46[4]\, \DATA_OUT_0_46[5]\, 
        \DATA_OUT_0_46[6]\, \DATA_OUT_0_46[7]\, 
        \DATA_OUT_0_46[8]\, \DATA_OUT_0_46[9]\, 
        \DATA_OUT_0_46[10]\, \DATA_OUT_0_46[11]\, 
        \DATA_OUT_0_46[12]\, \DATA_OUT_0_46[13]\, 
        \DATA_OUT_0_46[14]\, \DATA_OUT_0_46[15]\, 
        \DATA_OUT_0_46[16]\, \DATA_OUT_0_46[17]\, 
        \DATA_OUT_0_46[18]\, \DATA_OUT_0_46[19]\, 
        \DATA_OUT_0_46[20]\, \DATA_OUT_0_46[21]\, 
        \DATA_OUT_0_46[22]\, \DATA_OUT_0_46[23]\, 
        \DATA_OUT_0_46[24]\, \DATA_OUT_0_46[25]\, 
        \DATA_OUT_0_47[0]\, \DATA_OUT_0_47[1]\, 
        \DATA_OUT_0_47[2]\, \DATA_OUT_0_47[3]\, 
        \DATA_OUT_0_47[4]\, \DATA_OUT_0_47[5]\, 
        \DATA_OUT_0_47[6]\, \DATA_OUT_0_47[7]\, 
        \DATA_OUT_0_47[8]\, \DATA_OUT_0_47[9]\, 
        \DATA_OUT_0_47[10]\, \DATA_OUT_0_47[11]\, 
        \DATA_OUT_0_47[12]\, \DATA_OUT_0_47[13]\, 
        \DATA_OUT_0_47[14]\, \DATA_OUT_0_47[15]\, 
        \DATA_OUT_0_47[16]\, \DATA_OUT_0_47[17]\, 
        \DATA_OUT_0_47[18]\, \DATA_OUT_0_47[19]\, 
        \DATA_OUT_0_47[20]\, \DATA_OUT_0_47[21]\, 
        \DATA_OUT_0_47[22]\, \DATA_OUT_0_47[23]\, 
        \DATA_OUT_0_47[24]\, \DATA_OUT_0_47[25]\, 
        \DATA_OUT_0_48[0]\, \DATA_OUT_0_48[1]\, 
        \DATA_OUT_0_48[2]\, \DATA_OUT_0_48[3]\, 
        \DATA_OUT_0_48[4]\, \DATA_OUT_0_48[5]\, 
        \DATA_OUT_0_48[6]\, \DATA_OUT_0_48[7]\, 
        \DATA_OUT_0_48[8]\, \DATA_OUT_0_48[9]\, 
        \DATA_OUT_0_48[10]\, \DATA_OUT_0_48[11]\, 
        \DATA_OUT_0_48[12]\, \DATA_OUT_0_48[13]\, 
        \DATA_OUT_0_48[14]\, \DATA_OUT_0_48[15]\, 
        \DATA_OUT_0_48[16]\, \DATA_OUT_0_48[17]\, 
        \DATA_OUT_0_48[18]\, \DATA_OUT_0_48[19]\, 
        \DATA_OUT_0_48[20]\, \DATA_OUT_0_48[21]\, 
        \DATA_OUT_0_48[22]\, \DATA_OUT_0_48[23]\, 
        \DATA_OUT_0_48[24]\, \DATA_OUT_0_48[25]\, 
        \DATA_OUT_0_49[0]\, \DATA_OUT_0_49[1]\, 
        \DATA_OUT_0_49[2]\, \DATA_OUT_0_49[3]\, 
        \DATA_OUT_0_49[4]\, \DATA_OUT_0_49[5]\, 
        \DATA_OUT_0_49[6]\, \DATA_OUT_0_49[7]\, 
        \DATA_OUT_0_49[8]\, \DATA_OUT_0_49[9]\, 
        \DATA_OUT_0_49[10]\, \DATA_OUT_0_49[11]\, 
        \DATA_OUT_0_49[12]\, \DATA_OUT_0_49[13]\, 
        \DATA_OUT_0_49[14]\, \DATA_OUT_0_49[15]\, 
        \DATA_OUT_0_49[16]\, \DATA_OUT_0_49[17]\, 
        \DATA_OUT_0_49[18]\, \DATA_OUT_0_49[19]\, 
        \DATA_OUT_0_49[20]\, \DATA_OUT_0_49[21]\, 
        \DATA_OUT_0_49[22]\, \DATA_OUT_0_49[23]\, 
        \DATA_OUT_0_49[24]\, \DATA_OUT_0_49[25]\, 
        \DATA_OUT_0_50[0]\, \DATA_OUT_0_50[1]\, 
        \DATA_OUT_0_50[2]\, \DATA_OUT_0_50[3]\, 
        \DATA_OUT_0_50[4]\, \DATA_OUT_0_50[5]\, 
        \DATA_OUT_0_50[6]\, \DATA_OUT_0_50[7]\, 
        \DATA_OUT_0_50[8]\, \DATA_OUT_0_50[9]\, 
        \DATA_OUT_0_50[10]\, \DATA_OUT_0_50[11]\, 
        \DATA_OUT_0_50[12]\, \DATA_OUT_0_50[13]\, 
        \DATA_OUT_0_50[14]\, \DATA_OUT_0_50[15]\, 
        \DATA_OUT_0_50[16]\, \DATA_OUT_0_50[17]\, 
        \DATA_OUT_0_50[18]\, \DATA_OUT_0_50[19]\, 
        \DATA_OUT_0_50[20]\, \DATA_OUT_0_50[21]\, 
        \DATA_OUT_0_50[22]\, \DATA_OUT_0_50[23]\, 
        \DATA_OUT_0_50[24]\, \DATA_OUT_0_50[25]\, 
        \DATA_OUT_0_51[0]\, \DATA_OUT_0_51[1]\, 
        \DATA_OUT_0_51[2]\, \DATA_OUT_0_51[3]\, 
        \DATA_OUT_0_51[4]\, \DATA_OUT_0_51[5]\, 
        \DATA_OUT_0_51[6]\, \DATA_OUT_0_51[7]\, 
        \DATA_OUT_0_51[8]\, \DATA_OUT_0_51[9]\, 
        \DATA_OUT_0_51[10]\, \DATA_OUT_0_51[11]\, 
        \DATA_OUT_0_51[12]\, \DATA_OUT_0_51[13]\, 
        \DATA_OUT_0_51[14]\, \DATA_OUT_0_51[15]\, 
        \DATA_OUT_0_51[16]\, \DATA_OUT_0_51[17]\, 
        \DATA_OUT_0_51[18]\, \DATA_OUT_0_51[19]\, 
        \DATA_OUT_0_51[20]\, \DATA_OUT_0_51[21]\, 
        \DATA_OUT_0_51[22]\, \DATA_OUT_0_51[23]\, 
        \DATA_OUT_0_51[24]\, \DATA_OUT_0_51[25]\, 
        \DATA_OUT_1_0[0]\, \DATA_OUT_1_0[1]\, \DATA_OUT_1_0[2]\, 
        \DATA_OUT_1_0[3]\, \DATA_OUT_1_0[4]\, \DATA_OUT_1_0[5]\, 
        \DATA_OUT_1_0[6]\, \DATA_OUT_1_0[7]\, \DATA_OUT_1_0[8]\, 
        \DATA_OUT_1_0[9]\, \DATA_OUT_1_0[10]\, \DATA_OUT_1_0[11]\, 
        \DATA_OUT_1_0[12]\, \DATA_OUT_1_0[13]\, 
        \DATA_OUT_1_0[14]\, \DATA_OUT_1_0[15]\, 
        \DATA_OUT_1_0[16]\, \DATA_OUT_1_0[17]\, 
        \DATA_OUT_1_0[18]\, \DATA_OUT_1_0[19]\, 
        \DATA_OUT_1_0[20]\, \DATA_OUT_1_0[21]\, 
        \DATA_OUT_1_0[22]\, \DATA_OUT_1_0[23]\, 
        \DATA_OUT_1_0[24]\, \DATA_OUT_1_0[25]\, \DATA_OUT_1_1[0]\, 
        \DATA_OUT_1_1[1]\, \DATA_OUT_1_1[2]\, \DATA_OUT_1_1[3]\, 
        \DATA_OUT_1_1[4]\, \DATA_OUT_1_1[5]\, \DATA_OUT_1_1[6]\, 
        \DATA_OUT_1_1[7]\, \DATA_OUT_1_1[8]\, \DATA_OUT_1_1[9]\, 
        \DATA_OUT_1_1[10]\, \DATA_OUT_1_1[11]\, 
        \DATA_OUT_1_1[12]\, \DATA_OUT_1_1[13]\, 
        \DATA_OUT_1_1[14]\, \DATA_OUT_1_1[15]\, 
        \DATA_OUT_1_1[16]\, \DATA_OUT_1_1[17]\, 
        \DATA_OUT_1_1[18]\, \DATA_OUT_1_1[19]\, 
        \DATA_OUT_1_1[20]\, \DATA_OUT_1_1[21]\, 
        \DATA_OUT_1_1[22]\, \DATA_OUT_1_1[23]\, 
        \DATA_OUT_1_1[24]\, \DATA_OUT_1_1[25]\, \DATA_OUT_1_2[0]\, 
        \DATA_OUT_1_2[1]\, \DATA_OUT_1_2[2]\, \DATA_OUT_1_2[3]\, 
        \DATA_OUT_1_2[4]\, \DATA_OUT_1_2[5]\, \DATA_OUT_1_2[6]\, 
        \DATA_OUT_1_2[7]\, \DATA_OUT_1_2[8]\, \DATA_OUT_1_2[9]\, 
        \DATA_OUT_1_2[10]\, \DATA_OUT_1_2[11]\, 
        \DATA_OUT_1_2[12]\, \DATA_OUT_1_2[13]\, 
        \DATA_OUT_1_2[14]\, \DATA_OUT_1_2[15]\, 
        \DATA_OUT_1_2[16]\, \DATA_OUT_1_2[17]\, 
        \DATA_OUT_1_2[18]\, \DATA_OUT_1_2[19]\, 
        \DATA_OUT_1_2[20]\, \DATA_OUT_1_2[21]\, 
        \DATA_OUT_1_2[22]\, \DATA_OUT_1_2[23]\, 
        \DATA_OUT_1_2[24]\, \DATA_OUT_1_2[25]\, \DATA_OUT_1_3[0]\, 
        \DATA_OUT_1_3[1]\, \DATA_OUT_1_3[2]\, \DATA_OUT_1_3[3]\, 
        \DATA_OUT_1_3[4]\, \DATA_OUT_1_3[5]\, \DATA_OUT_1_3[6]\, 
        \DATA_OUT_1_3[7]\, \DATA_OUT_1_3[8]\, \DATA_OUT_1_3[9]\, 
        \DATA_OUT_1_3[10]\, \DATA_OUT_1_3[11]\, 
        \DATA_OUT_1_3[12]\, \DATA_OUT_1_3[13]\, 
        \DATA_OUT_1_3[14]\, \DATA_OUT_1_3[15]\, 
        \DATA_OUT_1_3[16]\, \DATA_OUT_1_3[17]\, 
        \DATA_OUT_1_3[18]\, \DATA_OUT_1_3[19]\, 
        \DATA_OUT_1_3[20]\, \DATA_OUT_1_3[21]\, 
        \DATA_OUT_1_3[22]\, \DATA_OUT_1_3[23]\, 
        \DATA_OUT_1_3[24]\, \DATA_OUT_1_3[25]\, \DATA_OUT_1_4[0]\, 
        \DATA_OUT_1_4[1]\, \DATA_OUT_1_4[2]\, \DATA_OUT_1_4[3]\, 
        \DATA_OUT_1_4[4]\, \DATA_OUT_1_4[5]\, \DATA_OUT_1_4[6]\, 
        \DATA_OUT_1_4[7]\, \DATA_OUT_1_4[8]\, \DATA_OUT_1_4[9]\, 
        \DATA_OUT_1_4[10]\, \DATA_OUT_1_4[11]\, 
        \DATA_OUT_1_4[12]\, \DATA_OUT_1_4[13]\, 
        \DATA_OUT_1_4[14]\, \DATA_OUT_1_4[15]\, 
        \DATA_OUT_1_4[16]\, \DATA_OUT_1_4[17]\, 
        \DATA_OUT_1_4[18]\, \DATA_OUT_1_4[19]\, 
        \DATA_OUT_1_4[20]\, \DATA_OUT_1_4[21]\, 
        \DATA_OUT_1_4[22]\, \DATA_OUT_1_4[23]\, 
        \DATA_OUT_1_4[24]\, \DATA_OUT_1_4[25]\, \DATA_OUT_1_5[0]\, 
        \DATA_OUT_1_5[1]\, \DATA_OUT_1_5[2]\, \DATA_OUT_1_5[3]\, 
        \DATA_OUT_1_5[4]\, \DATA_OUT_1_5[5]\, \DATA_OUT_1_5[6]\, 
        \DATA_OUT_1_5[7]\, \DATA_OUT_1_5[8]\, \DATA_OUT_1_5[9]\, 
        \DATA_OUT_1_5[10]\, \DATA_OUT_1_5[11]\, 
        \DATA_OUT_1_5[12]\, \DATA_OUT_1_5[13]\, 
        \DATA_OUT_1_5[14]\, \DATA_OUT_1_5[15]\, 
        \DATA_OUT_1_5[16]\, \DATA_OUT_1_5[17]\, 
        \DATA_OUT_1_5[18]\, \DATA_OUT_1_5[19]\, 
        \DATA_OUT_1_5[20]\, \DATA_OUT_1_5[21]\, 
        \DATA_OUT_1_5[22]\, \DATA_OUT_1_5[23]\, 
        \DATA_OUT_1_5[24]\, \DATA_OUT_1_5[25]\, \DATA_OUT_1_6[0]\, 
        \DATA_OUT_1_6[1]\, \DATA_OUT_1_6[2]\, \DATA_OUT_1_6[3]\, 
        \DATA_OUT_1_6[4]\, \DATA_OUT_1_6[5]\, \DATA_OUT_1_6[6]\, 
        \DATA_OUT_1_6[7]\, \DATA_OUT_1_6[8]\, \DATA_OUT_1_6[9]\, 
        \DATA_OUT_1_6[10]\, \DATA_OUT_1_6[11]\, 
        \DATA_OUT_1_6[12]\, \DATA_OUT_1_6[13]\, 
        \DATA_OUT_1_6[14]\, \DATA_OUT_1_6[15]\, 
        \DATA_OUT_1_6[16]\, \DATA_OUT_1_6[17]\, 
        \DATA_OUT_1_6[18]\, \DATA_OUT_1_6[19]\, 
        \DATA_OUT_1_6[20]\, \DATA_OUT_1_6[21]\, 
        \DATA_OUT_1_6[22]\, \DATA_OUT_1_6[23]\, 
        \DATA_OUT_1_6[24]\, \DATA_OUT_1_6[25]\, \DATA_OUT_1_7[0]\, 
        \DATA_OUT_1_7[1]\, \DATA_OUT_1_7[2]\, \DATA_OUT_1_7[3]\, 
        \DATA_OUT_1_7[4]\, \DATA_OUT_1_7[5]\, \DATA_OUT_1_7[6]\, 
        \DATA_OUT_1_7[7]\, \DATA_OUT_1_7[8]\, \DATA_OUT_1_7[9]\, 
        \DATA_OUT_1_7[10]\, \DATA_OUT_1_7[11]\, 
        \DATA_OUT_1_7[12]\, \DATA_OUT_1_7[13]\, 
        \DATA_OUT_1_7[14]\, \DATA_OUT_1_7[15]\, 
        \DATA_OUT_1_7[16]\, \DATA_OUT_1_7[17]\, 
        \DATA_OUT_1_7[18]\, \DATA_OUT_1_7[19]\, 
        \DATA_OUT_1_7[20]\, \DATA_OUT_1_7[21]\, 
        \DATA_OUT_1_7[22]\, \DATA_OUT_1_7[23]\, 
        \DATA_OUT_1_7[24]\, \DATA_OUT_1_7[25]\, \DATA_OUT_1_8[0]\, 
        \DATA_OUT_1_8[1]\, \DATA_OUT_1_8[2]\, \DATA_OUT_1_8[3]\, 
        \DATA_OUT_1_8[4]\, \DATA_OUT_1_8[5]\, \DATA_OUT_1_8[6]\, 
        \DATA_OUT_1_8[7]\, \DATA_OUT_1_8[8]\, \DATA_OUT_1_8[9]\, 
        \DATA_OUT_1_8[10]\, \DATA_OUT_1_8[11]\, 
        \DATA_OUT_1_8[12]\, \DATA_OUT_1_8[13]\, 
        \DATA_OUT_1_8[14]\, \DATA_OUT_1_8[15]\, 
        \DATA_OUT_1_8[16]\, \DATA_OUT_1_8[17]\, 
        \DATA_OUT_1_8[18]\, \DATA_OUT_1_8[19]\, 
        \DATA_OUT_1_8[20]\, \DATA_OUT_1_8[21]\, 
        \DATA_OUT_1_8[22]\, \DATA_OUT_1_8[23]\, 
        \DATA_OUT_1_8[24]\, \DATA_OUT_1_8[25]\, \DATA_OUT_1_9[0]\, 
        \DATA_OUT_1_9[1]\, \DATA_OUT_1_9[2]\, \DATA_OUT_1_9[3]\, 
        \DATA_OUT_1_9[4]\, \DATA_OUT_1_9[5]\, \DATA_OUT_1_9[6]\, 
        \DATA_OUT_1_9[7]\, \DATA_OUT_1_9[8]\, \DATA_OUT_1_9[9]\, 
        \DATA_OUT_1_9[10]\, \DATA_OUT_1_9[11]\, 
        \DATA_OUT_1_9[12]\, \DATA_OUT_1_9[13]\, 
        \DATA_OUT_1_9[14]\, \DATA_OUT_1_9[15]\, 
        \DATA_OUT_1_9[16]\, \DATA_OUT_1_9[17]\, 
        \DATA_OUT_1_9[18]\, \DATA_OUT_1_9[19]\, 
        \DATA_OUT_1_9[20]\, \DATA_OUT_1_9[21]\, 
        \DATA_OUT_1_9[22]\, \DATA_OUT_1_9[23]\, 
        \DATA_OUT_1_9[24]\, \DATA_OUT_1_9[25]\, 
        \DATA_OUT_1_10[0]\, \DATA_OUT_1_10[1]\, 
        \DATA_OUT_1_10[2]\, \DATA_OUT_1_10[3]\, 
        \DATA_OUT_1_10[4]\, \DATA_OUT_1_10[5]\, 
        \DATA_OUT_1_10[6]\, \DATA_OUT_1_10[7]\, 
        \DATA_OUT_1_10[8]\, \DATA_OUT_1_10[9]\, 
        \DATA_OUT_1_10[10]\, \DATA_OUT_1_10[11]\, 
        \DATA_OUT_1_10[12]\, \DATA_OUT_1_10[13]\, 
        \DATA_OUT_1_10[14]\, \DATA_OUT_1_10[15]\, 
        \DATA_OUT_1_10[16]\, \DATA_OUT_1_10[17]\, 
        \DATA_OUT_1_10[18]\, \DATA_OUT_1_10[19]\, 
        \DATA_OUT_1_10[20]\, \DATA_OUT_1_10[21]\, 
        \DATA_OUT_1_10[22]\, \DATA_OUT_1_10[23]\, 
        \DATA_OUT_1_10[24]\, \DATA_OUT_1_10[25]\, 
        \DATA_OUT_1_11[0]\, \DATA_OUT_1_11[1]\, 
        \DATA_OUT_1_11[2]\, \DATA_OUT_1_11[3]\, 
        \DATA_OUT_1_11[4]\, \DATA_OUT_1_11[5]\, 
        \DATA_OUT_1_11[6]\, \DATA_OUT_1_11[7]\, 
        \DATA_OUT_1_11[8]\, \DATA_OUT_1_11[9]\, 
        \DATA_OUT_1_11[10]\, \DATA_OUT_1_11[11]\, 
        \DATA_OUT_1_11[12]\, \DATA_OUT_1_11[13]\, 
        \DATA_OUT_1_11[14]\, \DATA_OUT_1_11[15]\, 
        \DATA_OUT_1_11[16]\, \DATA_OUT_1_11[17]\, 
        \DATA_OUT_1_11[18]\, \DATA_OUT_1_11[19]\, 
        \DATA_OUT_1_11[20]\, \DATA_OUT_1_11[21]\, 
        \DATA_OUT_1_11[22]\, \DATA_OUT_1_11[23]\, 
        \DATA_OUT_1_11[24]\, \DATA_OUT_1_11[25]\, 
        \DATA_OUT_1_12[0]\, \DATA_OUT_1_12[1]\, 
        \DATA_OUT_1_12[2]\, \DATA_OUT_1_12[3]\, 
        \DATA_OUT_1_12[4]\, \DATA_OUT_1_12[5]\, 
        \DATA_OUT_1_12[6]\, \DATA_OUT_1_12[7]\, 
        \DATA_OUT_1_12[8]\, \DATA_OUT_1_12[9]\, 
        \DATA_OUT_1_12[10]\, \DATA_OUT_1_12[11]\, 
        \DATA_OUT_1_12[12]\, \DATA_OUT_1_12[13]\, 
        \DATA_OUT_1_12[14]\, \DATA_OUT_1_12[15]\, 
        \DATA_OUT_1_12[16]\, \DATA_OUT_1_12[17]\, 
        \DATA_OUT_1_12[18]\, \DATA_OUT_1_12[19]\, 
        \DATA_OUT_1_12[20]\, \DATA_OUT_1_12[21]\, 
        \DATA_OUT_1_12[22]\, \DATA_OUT_1_12[23]\, 
        \DATA_OUT_1_12[24]\, \DATA_OUT_1_12[25]\, 
        \DATA_OUT_1_13[0]\, \DATA_OUT_1_13[1]\, 
        \DATA_OUT_1_13[2]\, \DATA_OUT_1_13[3]\, 
        \DATA_OUT_1_13[4]\, \DATA_OUT_1_13[5]\, 
        \DATA_OUT_1_13[6]\, \DATA_OUT_1_13[7]\, 
        \DATA_OUT_1_13[8]\, \DATA_OUT_1_13[9]\, 
        \DATA_OUT_1_13[10]\, \DATA_OUT_1_13[11]\, 
        \DATA_OUT_1_13[12]\, \DATA_OUT_1_13[13]\, 
        \DATA_OUT_1_13[14]\, \DATA_OUT_1_13[15]\, 
        \DATA_OUT_1_13[16]\, \DATA_OUT_1_13[17]\, 
        \DATA_OUT_1_13[18]\, \DATA_OUT_1_13[19]\, 
        \DATA_OUT_1_13[20]\, \DATA_OUT_1_13[21]\, 
        \DATA_OUT_1_13[22]\, \DATA_OUT_1_13[23]\, 
        \DATA_OUT_1_13[24]\, \DATA_OUT_1_13[25]\, 
        \DATA_OUT_1_14[0]\, \DATA_OUT_1_14[1]\, 
        \DATA_OUT_1_14[2]\, \DATA_OUT_1_14[3]\, 
        \DATA_OUT_1_14[4]\, \DATA_OUT_1_14[5]\, 
        \DATA_OUT_1_14[6]\, \DATA_OUT_1_14[7]\, 
        \DATA_OUT_1_14[8]\, \DATA_OUT_1_14[9]\, 
        \DATA_OUT_1_14[10]\, \DATA_OUT_1_14[11]\, 
        \DATA_OUT_1_14[12]\, \DATA_OUT_1_14[13]\, 
        \DATA_OUT_1_14[14]\, \DATA_OUT_1_14[15]\, 
        \DATA_OUT_1_14[16]\, \DATA_OUT_1_14[17]\, 
        \DATA_OUT_1_14[18]\, \DATA_OUT_1_14[19]\, 
        \DATA_OUT_1_14[20]\, \DATA_OUT_1_14[21]\, 
        \DATA_OUT_1_14[22]\, \DATA_OUT_1_14[23]\, 
        \DATA_OUT_1_14[24]\, \DATA_OUT_1_14[25]\, 
        \DATA_OUT_1_15[0]\, \DATA_OUT_1_15[1]\, 
        \DATA_OUT_1_15[2]\, \DATA_OUT_1_15[3]\, 
        \DATA_OUT_1_15[4]\, \DATA_OUT_1_15[5]\, 
        \DATA_OUT_1_15[6]\, \DATA_OUT_1_15[7]\, 
        \DATA_OUT_1_15[8]\, \DATA_OUT_1_15[9]\, 
        \DATA_OUT_1_15[10]\, \DATA_OUT_1_15[11]\, 
        \DATA_OUT_1_15[12]\, \DATA_OUT_1_15[13]\, 
        \DATA_OUT_1_15[14]\, \DATA_OUT_1_15[15]\, 
        \DATA_OUT_1_15[16]\, \DATA_OUT_1_15[17]\, 
        \DATA_OUT_1_15[18]\, \DATA_OUT_1_15[19]\, 
        \DATA_OUT_1_15[20]\, \DATA_OUT_1_15[21]\, 
        \DATA_OUT_1_15[22]\, \DATA_OUT_1_15[23]\, 
        \DATA_OUT_1_15[24]\, \DATA_OUT_1_15[25]\, 
        \DATA_OUT_1_16[0]\, \DATA_OUT_1_16[1]\, 
        \DATA_OUT_1_16[2]\, \DATA_OUT_1_16[3]\, 
        \DATA_OUT_1_16[4]\, \DATA_OUT_1_16[5]\, 
        \DATA_OUT_1_16[6]\, \DATA_OUT_1_16[7]\, 
        \DATA_OUT_1_16[8]\, \DATA_OUT_1_16[9]\, 
        \DATA_OUT_1_16[10]\, \DATA_OUT_1_16[11]\, 
        \DATA_OUT_1_16[12]\, \DATA_OUT_1_16[13]\, 
        \DATA_OUT_1_16[14]\, \DATA_OUT_1_16[15]\, 
        \DATA_OUT_1_16[16]\, \DATA_OUT_1_16[17]\, 
        \DATA_OUT_1_16[18]\, \DATA_OUT_1_16[19]\, 
        \DATA_OUT_1_16[20]\, \DATA_OUT_1_16[21]\, 
        \DATA_OUT_1_16[22]\, \DATA_OUT_1_16[23]\, 
        \DATA_OUT_1_16[24]\, \DATA_OUT_1_16[25]\, 
        \DATA_OUT_1_17[0]\, \DATA_OUT_1_17[1]\, 
        \DATA_OUT_1_17[2]\, \DATA_OUT_1_17[3]\, 
        \DATA_OUT_1_17[4]\, \DATA_OUT_1_17[5]\, 
        \DATA_OUT_1_17[6]\, \DATA_OUT_1_17[7]\, 
        \DATA_OUT_1_17[8]\, \DATA_OUT_1_17[9]\, 
        \DATA_OUT_1_17[10]\, \DATA_OUT_1_17[11]\, 
        \DATA_OUT_1_17[12]\, \DATA_OUT_1_17[13]\, 
        \DATA_OUT_1_17[14]\, \DATA_OUT_1_17[15]\, 
        \DATA_OUT_1_17[16]\, \DATA_OUT_1_17[17]\, 
        \DATA_OUT_1_17[18]\, \DATA_OUT_1_17[19]\, 
        \DATA_OUT_1_17[20]\, \DATA_OUT_1_17[21]\, 
        \DATA_OUT_1_17[22]\, \DATA_OUT_1_17[23]\, 
        \DATA_OUT_1_17[24]\, \DATA_OUT_1_17[25]\, 
        \DATA_OUT_1_18[0]\, \DATA_OUT_1_18[1]\, 
        \DATA_OUT_1_18[2]\, \DATA_OUT_1_18[3]\, 
        \DATA_OUT_1_18[4]\, \DATA_OUT_1_18[5]\, 
        \DATA_OUT_1_18[6]\, \DATA_OUT_1_18[7]\, 
        \DATA_OUT_1_18[8]\, \DATA_OUT_1_18[9]\, 
        \DATA_OUT_1_18[10]\, \DATA_OUT_1_18[11]\, 
        \DATA_OUT_1_18[12]\, \DATA_OUT_1_18[13]\, 
        \DATA_OUT_1_18[14]\, \DATA_OUT_1_18[15]\, 
        \DATA_OUT_1_18[16]\, \DATA_OUT_1_18[17]\, 
        \DATA_OUT_1_18[18]\, \DATA_OUT_1_18[19]\, 
        \DATA_OUT_1_18[20]\, \DATA_OUT_1_18[21]\, 
        \DATA_OUT_1_18[22]\, \DATA_OUT_1_18[23]\, 
        \DATA_OUT_1_18[24]\, \DATA_OUT_1_18[25]\, 
        \DATA_OUT_1_19[0]\, \DATA_OUT_1_19[1]\, 
        \DATA_OUT_1_19[2]\, \DATA_OUT_1_19[3]\, 
        \DATA_OUT_1_19[4]\, \DATA_OUT_1_19[5]\, 
        \DATA_OUT_1_19[6]\, \DATA_OUT_1_19[7]\, 
        \DATA_OUT_1_19[8]\, \DATA_OUT_1_19[9]\, 
        \DATA_OUT_1_19[10]\, \DATA_OUT_1_19[11]\, 
        \DATA_OUT_1_19[12]\, \DATA_OUT_1_19[13]\, 
        \DATA_OUT_1_19[14]\, \DATA_OUT_1_19[15]\, 
        \DATA_OUT_1_19[16]\, \DATA_OUT_1_19[17]\, 
        \DATA_OUT_1_19[18]\, \DATA_OUT_1_19[19]\, 
        \DATA_OUT_1_19[20]\, \DATA_OUT_1_19[21]\, 
        \DATA_OUT_1_19[22]\, \DATA_OUT_1_19[23]\, 
        \DATA_OUT_1_19[24]\, \DATA_OUT_1_19[25]\, 
        \DATA_OUT_1_20[0]\, \DATA_OUT_1_20[1]\, 
        \DATA_OUT_1_20[2]\, \DATA_OUT_1_20[3]\, 
        \DATA_OUT_1_20[4]\, \DATA_OUT_1_20[5]\, 
        \DATA_OUT_1_20[6]\, \DATA_OUT_1_20[7]\, 
        \DATA_OUT_1_20[8]\, \DATA_OUT_1_20[9]\, 
        \DATA_OUT_1_20[10]\, \DATA_OUT_1_20[11]\, 
        \DATA_OUT_1_20[12]\, \DATA_OUT_1_20[13]\, 
        \DATA_OUT_1_20[14]\, \DATA_OUT_1_20[15]\, 
        \DATA_OUT_1_20[16]\, \DATA_OUT_1_20[17]\, 
        \DATA_OUT_1_20[18]\, \DATA_OUT_1_20[19]\, 
        \DATA_OUT_1_20[20]\, \DATA_OUT_1_20[21]\, 
        \DATA_OUT_1_20[22]\, \DATA_OUT_1_20[23]\, 
        \DATA_OUT_1_20[24]\, \DATA_OUT_1_20[25]\, 
        \DATA_OUT_1_21[0]\, \DATA_OUT_1_21[1]\, 
        \DATA_OUT_1_21[2]\, \DATA_OUT_1_21[3]\, 
        \DATA_OUT_1_21[4]\, \DATA_OUT_1_21[5]\, 
        \DATA_OUT_1_21[6]\, \DATA_OUT_1_21[7]\, 
        \DATA_OUT_1_21[8]\, \DATA_OUT_1_21[9]\, 
        \DATA_OUT_1_21[10]\, \DATA_OUT_1_21[11]\, 
        \DATA_OUT_1_21[12]\, \DATA_OUT_1_21[13]\, 
        \DATA_OUT_1_21[14]\, \DATA_OUT_1_21[15]\, 
        \DATA_OUT_1_21[16]\, \DATA_OUT_1_21[17]\, 
        \DATA_OUT_1_21[18]\, \DATA_OUT_1_21[19]\, 
        \DATA_OUT_1_21[20]\, \DATA_OUT_1_21[21]\, 
        \DATA_OUT_1_21[22]\, \DATA_OUT_1_21[23]\, 
        \DATA_OUT_1_21[24]\, \DATA_OUT_1_21[25]\, 
        \DATA_OUT_1_22[0]\, \DATA_OUT_1_22[1]\, 
        \DATA_OUT_1_22[2]\, \DATA_OUT_1_22[3]\, 
        \DATA_OUT_1_22[4]\, \DATA_OUT_1_22[5]\, 
        \DATA_OUT_1_22[6]\, \DATA_OUT_1_22[7]\, 
        \DATA_OUT_1_22[8]\, \DATA_OUT_1_22[9]\, 
        \DATA_OUT_1_22[10]\, \DATA_OUT_1_22[11]\, 
        \DATA_OUT_1_22[12]\, \DATA_OUT_1_22[13]\, 
        \DATA_OUT_1_22[14]\, \DATA_OUT_1_22[15]\, 
        \DATA_OUT_1_22[16]\, \DATA_OUT_1_22[17]\, 
        \DATA_OUT_1_22[18]\, \DATA_OUT_1_22[19]\, 
        \DATA_OUT_1_22[20]\, \DATA_OUT_1_22[21]\, 
        \DATA_OUT_1_22[22]\, \DATA_OUT_1_22[23]\, 
        \DATA_OUT_1_22[24]\, \DATA_OUT_1_22[25]\, 
        \DATA_OUT_1_23[0]\, \DATA_OUT_1_23[1]\, 
        \DATA_OUT_1_23[2]\, \DATA_OUT_1_23[3]\, 
        \DATA_OUT_1_23[4]\, \DATA_OUT_1_23[5]\, 
        \DATA_OUT_1_23[6]\, \DATA_OUT_1_23[7]\, 
        \DATA_OUT_1_23[8]\, \DATA_OUT_1_23[9]\, 
        \DATA_OUT_1_23[10]\, \DATA_OUT_1_23[11]\, 
        \DATA_OUT_1_23[12]\, \DATA_OUT_1_23[13]\, 
        \DATA_OUT_1_23[14]\, \DATA_OUT_1_23[15]\, 
        \DATA_OUT_1_23[16]\, \DATA_OUT_1_23[17]\, 
        \DATA_OUT_1_23[18]\, \DATA_OUT_1_23[19]\, 
        \DATA_OUT_1_23[20]\, \DATA_OUT_1_23[21]\, 
        \DATA_OUT_1_23[22]\, \DATA_OUT_1_23[23]\, 
        \DATA_OUT_1_23[24]\, \DATA_OUT_1_23[25]\, 
        \DATA_OUT_1_24[0]\, \DATA_OUT_1_24[1]\, 
        \DATA_OUT_1_24[2]\, \DATA_OUT_1_24[3]\, 
        \DATA_OUT_1_24[4]\, \DATA_OUT_1_24[5]\, 
        \DATA_OUT_1_24[6]\, \DATA_OUT_1_24[7]\, 
        \DATA_OUT_1_24[8]\, \DATA_OUT_1_24[9]\, 
        \DATA_OUT_1_24[10]\, \DATA_OUT_1_24[11]\, 
        \DATA_OUT_1_24[12]\, \DATA_OUT_1_24[13]\, 
        \DATA_OUT_1_24[14]\, \DATA_OUT_1_24[15]\, 
        \DATA_OUT_1_24[16]\, \DATA_OUT_1_24[17]\, 
        \DATA_OUT_1_24[18]\, \DATA_OUT_1_24[19]\, 
        \DATA_OUT_1_24[20]\, \DATA_OUT_1_24[21]\, 
        \DATA_OUT_1_24[22]\, \DATA_OUT_1_24[23]\, 
        \DATA_OUT_1_24[24]\, \DATA_OUT_1_24[25]\, 
        \DATA_OUT_1_25[0]\, \DATA_OUT_1_25[1]\, 
        \DATA_OUT_1_25[2]\, \DATA_OUT_1_25[3]\, 
        \DATA_OUT_1_25[4]\, \DATA_OUT_1_25[5]\, 
        \DATA_OUT_1_25[6]\, \DATA_OUT_1_25[7]\, 
        \DATA_OUT_1_25[8]\, \DATA_OUT_1_25[9]\, 
        \DATA_OUT_1_25[10]\, \DATA_OUT_1_25[11]\, 
        \DATA_OUT_1_25[12]\, \DATA_OUT_1_25[13]\, 
        \DATA_OUT_1_25[14]\, \DATA_OUT_1_25[15]\, 
        \DATA_OUT_1_25[16]\, \DATA_OUT_1_25[17]\, 
        \DATA_OUT_1_25[18]\, \DATA_OUT_1_25[19]\, 
        \DATA_OUT_1_25[20]\, \DATA_OUT_1_25[21]\, 
        \DATA_OUT_1_25[22]\, \DATA_OUT_1_25[23]\, 
        \DATA_OUT_1_25[24]\, \DATA_OUT_1_25[25]\, 
        \DATA_OUT_1_26[0]\, \DATA_OUT_1_26[1]\, 
        \DATA_OUT_1_26[2]\, \DATA_OUT_1_26[3]\, 
        \DATA_OUT_1_26[4]\, \DATA_OUT_1_26[5]\, 
        \DATA_OUT_1_26[6]\, \DATA_OUT_1_26[7]\, 
        \DATA_OUT_1_26[8]\, \DATA_OUT_1_26[9]\, 
        \DATA_OUT_1_26[10]\, \DATA_OUT_1_26[11]\, 
        \DATA_OUT_1_26[12]\, \DATA_OUT_1_26[13]\, 
        \DATA_OUT_1_26[14]\, \DATA_OUT_1_26[15]\, 
        \DATA_OUT_1_26[16]\, \DATA_OUT_1_26[17]\, 
        \DATA_OUT_1_26[18]\, \DATA_OUT_1_26[19]\, 
        \DATA_OUT_1_26[20]\, \DATA_OUT_1_26[21]\, 
        \DATA_OUT_1_26[22]\, \DATA_OUT_1_26[23]\, 
        \DATA_OUT_1_26[24]\, \DATA_OUT_1_26[25]\, 
        \DATA_OUT_1_27[0]\, \DATA_OUT_1_27[1]\, 
        \DATA_OUT_1_27[2]\, \DATA_OUT_1_27[3]\, 
        \DATA_OUT_1_27[4]\, \DATA_OUT_1_27[5]\, 
        \DATA_OUT_1_27[6]\, \DATA_OUT_1_27[7]\, 
        \DATA_OUT_1_27[8]\, \DATA_OUT_1_27[9]\, 
        \DATA_OUT_1_27[10]\, \DATA_OUT_1_27[11]\, 
        \DATA_OUT_1_27[12]\, \DATA_OUT_1_27[13]\, 
        \DATA_OUT_1_27[14]\, \DATA_OUT_1_27[15]\, 
        \DATA_OUT_1_27[16]\, \DATA_OUT_1_27[17]\, 
        \DATA_OUT_1_27[18]\, \DATA_OUT_1_27[19]\, 
        \DATA_OUT_1_27[20]\, \DATA_OUT_1_27[21]\, 
        \DATA_OUT_1_27[22]\, \DATA_OUT_1_27[23]\, 
        \DATA_OUT_1_27[24]\, \DATA_OUT_1_27[25]\, 
        \DATA_OUT_1_28[0]\, \DATA_OUT_1_28[1]\, 
        \DATA_OUT_1_28[2]\, \DATA_OUT_1_28[3]\, 
        \DATA_OUT_1_28[4]\, \DATA_OUT_1_28[5]\, 
        \DATA_OUT_1_28[6]\, \DATA_OUT_1_28[7]\, 
        \DATA_OUT_1_28[8]\, \DATA_OUT_1_28[9]\, 
        \DATA_OUT_1_28[10]\, \DATA_OUT_1_28[11]\, 
        \DATA_OUT_1_28[12]\, \DATA_OUT_1_28[13]\, 
        \DATA_OUT_1_28[14]\, \DATA_OUT_1_28[15]\, 
        \DATA_OUT_1_28[16]\, \DATA_OUT_1_28[17]\, 
        \DATA_OUT_1_28[18]\, \DATA_OUT_1_28[19]\, 
        \DATA_OUT_1_28[20]\, \DATA_OUT_1_28[21]\, 
        \DATA_OUT_1_28[22]\, \DATA_OUT_1_28[23]\, 
        \DATA_OUT_1_28[24]\, \DATA_OUT_1_28[25]\, 
        \DATA_OUT_1_29[0]\, \DATA_OUT_1_29[1]\, 
        \DATA_OUT_1_29[2]\, \DATA_OUT_1_29[3]\, 
        \DATA_OUT_1_29[4]\, \DATA_OUT_1_29[5]\, 
        \DATA_OUT_1_29[6]\, \DATA_OUT_1_29[7]\, 
        \DATA_OUT_1_29[8]\, \DATA_OUT_1_29[9]\, 
        \DATA_OUT_1_29[10]\, \DATA_OUT_1_29[11]\, 
        \DATA_OUT_1_29[12]\, \DATA_OUT_1_29[13]\, 
        \DATA_OUT_1_29[14]\, \DATA_OUT_1_29[15]\, 
        \DATA_OUT_1_29[16]\, \DATA_OUT_1_29[17]\, 
        \DATA_OUT_1_29[18]\, \DATA_OUT_1_29[19]\, 
        \DATA_OUT_1_29[20]\, \DATA_OUT_1_29[21]\, 
        \DATA_OUT_1_29[22]\, \DATA_OUT_1_29[23]\, 
        \DATA_OUT_1_29[24]\, \DATA_OUT_1_29[25]\, 
        \DATA_OUT_1_30[0]\, \DATA_OUT_1_30[1]\, 
        \DATA_OUT_1_30[2]\, \DATA_OUT_1_30[3]\, 
        \DATA_OUT_1_30[4]\, \DATA_OUT_1_30[5]\, 
        \DATA_OUT_1_30[6]\, \DATA_OUT_1_30[7]\, 
        \DATA_OUT_1_30[8]\, \DATA_OUT_1_30[9]\, 
        \DATA_OUT_1_30[10]\, \DATA_OUT_1_30[11]\, 
        \DATA_OUT_1_30[12]\, \DATA_OUT_1_30[13]\, 
        \DATA_OUT_1_30[14]\, \DATA_OUT_1_30[15]\, 
        \DATA_OUT_1_30[16]\, \DATA_OUT_1_30[17]\, 
        \DATA_OUT_1_30[18]\, \DATA_OUT_1_30[19]\, 
        \DATA_OUT_1_30[20]\, \DATA_OUT_1_30[21]\, 
        \DATA_OUT_1_30[22]\, \DATA_OUT_1_30[23]\, 
        \DATA_OUT_1_30[24]\, \DATA_OUT_1_30[25]\, 
        \DATA_OUT_1_31[0]\, \DATA_OUT_1_31[1]\, 
        \DATA_OUT_1_31[2]\, \DATA_OUT_1_31[3]\, 
        \DATA_OUT_1_31[4]\, \DATA_OUT_1_31[5]\, 
        \DATA_OUT_1_31[6]\, \DATA_OUT_1_31[7]\, 
        \DATA_OUT_1_31[8]\, \DATA_OUT_1_31[9]\, 
        \DATA_OUT_1_31[10]\, \DATA_OUT_1_31[11]\, 
        \DATA_OUT_1_31[12]\, \DATA_OUT_1_31[13]\, 
        \DATA_OUT_1_31[14]\, \DATA_OUT_1_31[15]\, 
        \DATA_OUT_1_31[16]\, \DATA_OUT_1_31[17]\, 
        \DATA_OUT_1_31[18]\, \DATA_OUT_1_31[19]\, 
        \DATA_OUT_1_31[20]\, \DATA_OUT_1_31[21]\, 
        \DATA_OUT_1_31[22]\, \DATA_OUT_1_31[23]\, 
        \DATA_OUT_1_31[24]\, \DATA_OUT_1_31[25]\, 
        \DATA_OUT_1_32[0]\, \DATA_OUT_1_32[1]\, 
        \DATA_OUT_1_32[2]\, \DATA_OUT_1_32[3]\, 
        \DATA_OUT_1_32[4]\, \DATA_OUT_1_32[5]\, 
        \DATA_OUT_1_32[6]\, \DATA_OUT_1_32[7]\, 
        \DATA_OUT_1_32[8]\, \DATA_OUT_1_32[9]\, 
        \DATA_OUT_1_32[10]\, \DATA_OUT_1_32[11]\, 
        \DATA_OUT_1_32[12]\, \DATA_OUT_1_32[13]\, 
        \DATA_OUT_1_32[14]\, \DATA_OUT_1_32[15]\, 
        \DATA_OUT_1_32[16]\, \DATA_OUT_1_32[17]\, 
        \DATA_OUT_1_32[18]\, \DATA_OUT_1_32[19]\, 
        \DATA_OUT_1_32[20]\, \DATA_OUT_1_32[21]\, 
        \DATA_OUT_1_32[22]\, \DATA_OUT_1_32[23]\, 
        \DATA_OUT_1_32[24]\, \DATA_OUT_1_32[25]\, 
        \DATA_OUT_1_33[0]\, \DATA_OUT_1_33[1]\, 
        \DATA_OUT_1_33[2]\, \DATA_OUT_1_33[3]\, 
        \DATA_OUT_1_33[4]\, \DATA_OUT_1_33[5]\, 
        \DATA_OUT_1_33[6]\, \DATA_OUT_1_33[7]\, 
        \DATA_OUT_1_33[8]\, \DATA_OUT_1_33[9]\, 
        \DATA_OUT_1_33[10]\, \DATA_OUT_1_33[11]\, 
        \DATA_OUT_1_33[12]\, \DATA_OUT_1_33[13]\, 
        \DATA_OUT_1_33[14]\, \DATA_OUT_1_33[15]\, 
        \DATA_OUT_1_33[16]\, \DATA_OUT_1_33[17]\, 
        \DATA_OUT_1_33[18]\, \DATA_OUT_1_33[19]\, 
        \DATA_OUT_1_33[20]\, \DATA_OUT_1_33[21]\, 
        \DATA_OUT_1_33[22]\, \DATA_OUT_1_33[23]\, 
        \DATA_OUT_1_33[24]\, \DATA_OUT_1_33[25]\, 
        \DATA_OUT_1_34[0]\, \DATA_OUT_1_34[1]\, 
        \DATA_OUT_1_34[2]\, \DATA_OUT_1_34[3]\, 
        \DATA_OUT_1_34[4]\, \DATA_OUT_1_34[5]\, 
        \DATA_OUT_1_34[6]\, \DATA_OUT_1_34[7]\, 
        \DATA_OUT_1_34[8]\, \DATA_OUT_1_34[9]\, 
        \DATA_OUT_1_34[10]\, \DATA_OUT_1_34[11]\, 
        \DATA_OUT_1_34[12]\, \DATA_OUT_1_34[13]\, 
        \DATA_OUT_1_34[14]\, \DATA_OUT_1_34[15]\, 
        \DATA_OUT_1_34[16]\, \DATA_OUT_1_34[17]\, 
        \DATA_OUT_1_34[18]\, \DATA_OUT_1_34[19]\, 
        \DATA_OUT_1_34[20]\, \DATA_OUT_1_34[21]\, 
        \DATA_OUT_1_34[22]\, \DATA_OUT_1_34[23]\, 
        \DATA_OUT_1_34[24]\, \DATA_OUT_1_34[25]\, 
        \DATA_OUT_1_35[0]\, \DATA_OUT_1_35[1]\, 
        \DATA_OUT_1_35[2]\, \DATA_OUT_1_35[3]\, 
        \DATA_OUT_1_35[4]\, \DATA_OUT_1_35[5]\, 
        \DATA_OUT_1_35[6]\, \DATA_OUT_1_35[7]\, 
        \DATA_OUT_1_35[8]\, \DATA_OUT_1_35[9]\, 
        \DATA_OUT_1_35[10]\, \DATA_OUT_1_35[11]\, 
        \DATA_OUT_1_35[12]\, \DATA_OUT_1_35[13]\, 
        \DATA_OUT_1_35[14]\, \DATA_OUT_1_35[15]\, 
        \DATA_OUT_1_35[16]\, \DATA_OUT_1_35[17]\, 
        \DATA_OUT_1_35[18]\, \DATA_OUT_1_35[19]\, 
        \DATA_OUT_1_35[20]\, \DATA_OUT_1_35[21]\, 
        \DATA_OUT_1_35[22]\, \DATA_OUT_1_35[23]\, 
        \DATA_OUT_1_35[24]\, \DATA_OUT_1_35[25]\, 
        \DATA_OUT_1_36[0]\, \DATA_OUT_1_36[1]\, 
        \DATA_OUT_1_36[2]\, \DATA_OUT_1_36[3]\, 
        \DATA_OUT_1_36[4]\, \DATA_OUT_1_36[5]\, 
        \DATA_OUT_1_36[6]\, \DATA_OUT_1_36[7]\, 
        \DATA_OUT_1_36[8]\, \DATA_OUT_1_36[9]\, 
        \DATA_OUT_1_36[10]\, \DATA_OUT_1_36[11]\, 
        \DATA_OUT_1_36[12]\, \DATA_OUT_1_36[13]\, 
        \DATA_OUT_1_36[14]\, \DATA_OUT_1_36[15]\, 
        \DATA_OUT_1_36[16]\, \DATA_OUT_1_36[17]\, 
        \DATA_OUT_1_36[18]\, \DATA_OUT_1_36[19]\, 
        \DATA_OUT_1_36[20]\, \DATA_OUT_1_36[21]\, 
        \DATA_OUT_1_36[22]\, \DATA_OUT_1_36[23]\, 
        \DATA_OUT_1_36[24]\, \DATA_OUT_1_36[25]\, 
        \DATA_OUT_1_37[0]\, \DATA_OUT_1_37[1]\, 
        \DATA_OUT_1_37[2]\, \DATA_OUT_1_37[3]\, 
        \DATA_OUT_1_37[4]\, \DATA_OUT_1_37[5]\, 
        \DATA_OUT_1_37[6]\, \DATA_OUT_1_37[7]\, 
        \DATA_OUT_1_37[8]\, \DATA_OUT_1_37[9]\, 
        \DATA_OUT_1_37[10]\, \DATA_OUT_1_37[11]\, 
        \DATA_OUT_1_37[12]\, \DATA_OUT_1_37[13]\, 
        \DATA_OUT_1_37[14]\, \DATA_OUT_1_37[15]\, 
        \DATA_OUT_1_37[16]\, \DATA_OUT_1_37[17]\, 
        \DATA_OUT_1_37[18]\, \DATA_OUT_1_37[19]\, 
        \DATA_OUT_1_37[20]\, \DATA_OUT_1_37[21]\, 
        \DATA_OUT_1_37[22]\, \DATA_OUT_1_37[23]\, 
        \DATA_OUT_1_37[24]\, \DATA_OUT_1_37[25]\, 
        \DATA_OUT_1_38[0]\, \DATA_OUT_1_38[1]\, 
        \DATA_OUT_1_38[2]\, \DATA_OUT_1_38[3]\, 
        \DATA_OUT_1_38[4]\, \DATA_OUT_1_38[5]\, 
        \DATA_OUT_1_38[6]\, \DATA_OUT_1_38[7]\, 
        \DATA_OUT_1_38[8]\, \DATA_OUT_1_38[9]\, 
        \DATA_OUT_1_38[10]\, \DATA_OUT_1_38[11]\, 
        \DATA_OUT_1_38[12]\, \DATA_OUT_1_38[13]\, 
        \DATA_OUT_1_38[14]\, \DATA_OUT_1_38[15]\, 
        \DATA_OUT_1_38[16]\, \DATA_OUT_1_38[17]\, 
        \DATA_OUT_1_38[18]\, \DATA_OUT_1_38[19]\, 
        \DATA_OUT_1_38[20]\, \DATA_OUT_1_38[21]\, 
        \DATA_OUT_1_38[22]\, \DATA_OUT_1_38[23]\, 
        \DATA_OUT_1_38[24]\, \DATA_OUT_1_38[25]\, 
        \DATA_OUT_1_39[0]\, \DATA_OUT_1_39[1]\, 
        \DATA_OUT_1_39[2]\, \DATA_OUT_1_39[3]\, 
        \DATA_OUT_1_39[4]\, \DATA_OUT_1_39[5]\, 
        \DATA_OUT_1_39[6]\, \DATA_OUT_1_39[7]\, 
        \DATA_OUT_1_39[8]\, \DATA_OUT_1_39[9]\, 
        \DATA_OUT_1_39[10]\, \DATA_OUT_1_39[11]\, 
        \DATA_OUT_1_39[12]\, \DATA_OUT_1_39[13]\, 
        \DATA_OUT_1_39[14]\, \DATA_OUT_1_39[15]\, 
        \DATA_OUT_1_39[16]\, \DATA_OUT_1_39[17]\, 
        \DATA_OUT_1_39[18]\, \DATA_OUT_1_39[19]\, 
        \DATA_OUT_1_39[20]\, \DATA_OUT_1_39[21]\, 
        \DATA_OUT_1_39[22]\, \DATA_OUT_1_39[23]\, 
        \DATA_OUT_1_39[24]\, \DATA_OUT_1_39[25]\, 
        \DATA_OUT_1_40[0]\, \DATA_OUT_1_40[1]\, 
        \DATA_OUT_1_40[2]\, \DATA_OUT_1_40[3]\, 
        \DATA_OUT_1_40[4]\, \DATA_OUT_1_40[5]\, 
        \DATA_OUT_1_40[6]\, \DATA_OUT_1_40[7]\, 
        \DATA_OUT_1_40[8]\, \DATA_OUT_1_40[9]\, 
        \DATA_OUT_1_40[10]\, \DATA_OUT_1_40[11]\, 
        \DATA_OUT_1_40[12]\, \DATA_OUT_1_40[13]\, 
        \DATA_OUT_1_40[14]\, \DATA_OUT_1_40[15]\, 
        \DATA_OUT_1_40[16]\, \DATA_OUT_1_40[17]\, 
        \DATA_OUT_1_40[18]\, \DATA_OUT_1_40[19]\, 
        \DATA_OUT_1_40[20]\, \DATA_OUT_1_40[21]\, 
        \DATA_OUT_1_40[22]\, \DATA_OUT_1_40[23]\, 
        \DATA_OUT_1_40[24]\, \DATA_OUT_1_40[25]\, 
        \DATA_OUT_1_41[0]\, \DATA_OUT_1_41[1]\, 
        \DATA_OUT_1_41[2]\, \DATA_OUT_1_41[3]\, 
        \DATA_OUT_1_41[4]\, \DATA_OUT_1_41[5]\, 
        \DATA_OUT_1_41[6]\, \DATA_OUT_1_41[7]\, 
        \DATA_OUT_1_41[8]\, \DATA_OUT_1_41[9]\, 
        \DATA_OUT_1_41[10]\, \DATA_OUT_1_41[11]\, 
        \DATA_OUT_1_41[12]\, \DATA_OUT_1_41[13]\, 
        \DATA_OUT_1_41[14]\, \DATA_OUT_1_41[15]\, 
        \DATA_OUT_1_41[16]\, \DATA_OUT_1_41[17]\, 
        \DATA_OUT_1_41[18]\, \DATA_OUT_1_41[19]\, 
        \DATA_OUT_1_41[20]\, \DATA_OUT_1_41[21]\, 
        \DATA_OUT_1_41[22]\, \DATA_OUT_1_41[23]\, 
        \DATA_OUT_1_41[24]\, \DATA_OUT_1_41[25]\, 
        \DATA_OUT_1_42[0]\, \DATA_OUT_1_42[1]\, 
        \DATA_OUT_1_42[2]\, \DATA_OUT_1_42[3]\, 
        \DATA_OUT_1_42[4]\, \DATA_OUT_1_42[5]\, 
        \DATA_OUT_1_42[6]\, \DATA_OUT_1_42[7]\, 
        \DATA_OUT_1_42[8]\, \DATA_OUT_1_42[9]\, 
        \DATA_OUT_1_42[10]\, \DATA_OUT_1_42[11]\, 
        \DATA_OUT_1_42[12]\, \DATA_OUT_1_42[13]\, 
        \DATA_OUT_1_42[14]\, \DATA_OUT_1_42[15]\, 
        \DATA_OUT_1_42[16]\, \DATA_OUT_1_42[17]\, 
        \DATA_OUT_1_42[18]\, \DATA_OUT_1_42[19]\, 
        \DATA_OUT_1_42[20]\, \DATA_OUT_1_42[21]\, 
        \DATA_OUT_1_42[22]\, \DATA_OUT_1_42[23]\, 
        \DATA_OUT_1_42[24]\, \DATA_OUT_1_42[25]\, 
        \DATA_OUT_1_43[0]\, \DATA_OUT_1_43[1]\, 
        \DATA_OUT_1_43[2]\, \DATA_OUT_1_43[3]\, 
        \DATA_OUT_1_43[4]\, \DATA_OUT_1_43[5]\, 
        \DATA_OUT_1_43[6]\, \DATA_OUT_1_43[7]\, 
        \DATA_OUT_1_43[8]\, \DATA_OUT_1_43[9]\, 
        \DATA_OUT_1_43[10]\, \DATA_OUT_1_43[11]\, 
        \DATA_OUT_1_43[12]\, \DATA_OUT_1_43[13]\, 
        \DATA_OUT_1_43[14]\, \DATA_OUT_1_43[15]\, 
        \DATA_OUT_1_43[16]\, \DATA_OUT_1_43[17]\, 
        \DATA_OUT_1_43[18]\, \DATA_OUT_1_43[19]\, 
        \DATA_OUT_1_43[20]\, \DATA_OUT_1_43[21]\, 
        \DATA_OUT_1_43[22]\, \DATA_OUT_1_43[23]\, 
        \DATA_OUT_1_43[24]\, \DATA_OUT_1_43[25]\, 
        \DATA_OUT_1_44[0]\, \DATA_OUT_1_44[1]\, 
        \DATA_OUT_1_44[2]\, \DATA_OUT_1_44[3]\, 
        \DATA_OUT_1_44[4]\, \DATA_OUT_1_44[5]\, 
        \DATA_OUT_1_44[6]\, \DATA_OUT_1_44[7]\, 
        \DATA_OUT_1_44[8]\, \DATA_OUT_1_44[9]\, 
        \DATA_OUT_1_44[10]\, \DATA_OUT_1_44[11]\, 
        \DATA_OUT_1_44[12]\, \DATA_OUT_1_44[13]\, 
        \DATA_OUT_1_44[14]\, \DATA_OUT_1_44[15]\, 
        \DATA_OUT_1_44[16]\, \DATA_OUT_1_44[17]\, 
        \DATA_OUT_1_44[18]\, \DATA_OUT_1_44[19]\, 
        \DATA_OUT_1_44[20]\, \DATA_OUT_1_44[21]\, 
        \DATA_OUT_1_44[22]\, \DATA_OUT_1_44[23]\, 
        \DATA_OUT_1_44[24]\, \DATA_OUT_1_44[25]\, 
        \DATA_OUT_1_45[0]\, \DATA_OUT_1_45[1]\, 
        \DATA_OUT_1_45[2]\, \DATA_OUT_1_45[3]\, 
        \DATA_OUT_1_45[4]\, \DATA_OUT_1_45[5]\, 
        \DATA_OUT_1_45[6]\, \DATA_OUT_1_45[7]\, 
        \DATA_OUT_1_45[8]\, \DATA_OUT_1_45[9]\, 
        \DATA_OUT_1_45[10]\, \DATA_OUT_1_45[11]\, 
        \DATA_OUT_1_45[12]\, \DATA_OUT_1_45[13]\, 
        \DATA_OUT_1_45[14]\, \DATA_OUT_1_45[15]\, 
        \DATA_OUT_1_45[16]\, \DATA_OUT_1_45[17]\, 
        \DATA_OUT_1_45[18]\, \DATA_OUT_1_45[19]\, 
        \DATA_OUT_1_45[20]\, \DATA_OUT_1_45[21]\, 
        \DATA_OUT_1_45[22]\, \DATA_OUT_1_45[23]\, 
        \DATA_OUT_1_45[24]\, \DATA_OUT_1_45[25]\, 
        \DATA_OUT_1_46[0]\, \DATA_OUT_1_46[1]\, 
        \DATA_OUT_1_46[2]\, \DATA_OUT_1_46[3]\, 
        \DATA_OUT_1_46[4]\, \DATA_OUT_1_46[5]\, 
        \DATA_OUT_1_46[6]\, \DATA_OUT_1_46[7]\, 
        \DATA_OUT_1_46[8]\, \DATA_OUT_1_46[9]\, 
        \DATA_OUT_1_46[10]\, \DATA_OUT_1_46[11]\, 
        \DATA_OUT_1_46[12]\, \DATA_OUT_1_46[13]\, 
        \DATA_OUT_1_46[14]\, \DATA_OUT_1_46[15]\, 
        \DATA_OUT_1_46[16]\, \DATA_OUT_1_46[17]\, 
        \DATA_OUT_1_46[18]\, \DATA_OUT_1_46[19]\, 
        \DATA_OUT_1_46[20]\, \DATA_OUT_1_46[21]\, 
        \DATA_OUT_1_46[22]\, \DATA_OUT_1_46[23]\, 
        \DATA_OUT_1_46[24]\, \DATA_OUT_1_46[25]\, 
        \DATA_OUT_1_47[0]\, \DATA_OUT_1_47[1]\, 
        \DATA_OUT_1_47[2]\, \DATA_OUT_1_47[3]\, 
        \DATA_OUT_1_47[4]\, \DATA_OUT_1_47[5]\, 
        \DATA_OUT_1_47[6]\, \DATA_OUT_1_47[7]\, 
        \DATA_OUT_1_47[8]\, \DATA_OUT_1_47[9]\, 
        \DATA_OUT_1_47[10]\, \DATA_OUT_1_47[11]\, 
        \DATA_OUT_1_47[12]\, \DATA_OUT_1_47[13]\, 
        \DATA_OUT_1_47[14]\, \DATA_OUT_1_47[15]\, 
        \DATA_OUT_1_47[16]\, \DATA_OUT_1_47[17]\, 
        \DATA_OUT_1_47[18]\, \DATA_OUT_1_47[19]\, 
        \DATA_OUT_1_47[20]\, \DATA_OUT_1_47[21]\, 
        \DATA_OUT_1_47[22]\, \DATA_OUT_1_47[23]\, 
        \DATA_OUT_1_47[24]\, \DATA_OUT_1_47[25]\, 
        \DATA_OUT_1_48[0]\, \DATA_OUT_1_48[1]\, 
        \DATA_OUT_1_48[2]\, \DATA_OUT_1_48[3]\, 
        \DATA_OUT_1_48[4]\, \DATA_OUT_1_48[5]\, 
        \DATA_OUT_1_48[6]\, \DATA_OUT_1_48[7]\, 
        \DATA_OUT_1_48[8]\, \DATA_OUT_1_48[9]\, 
        \DATA_OUT_1_48[10]\, \DATA_OUT_1_48[11]\, 
        \DATA_OUT_1_48[12]\, \DATA_OUT_1_48[13]\, 
        \DATA_OUT_1_48[14]\, \DATA_OUT_1_48[15]\, 
        \DATA_OUT_1_48[16]\, \DATA_OUT_1_48[17]\, 
        \DATA_OUT_1_48[18]\, \DATA_OUT_1_48[19]\, 
        \DATA_OUT_1_48[20]\, \DATA_OUT_1_48[21]\, 
        \DATA_OUT_1_48[22]\, \DATA_OUT_1_48[23]\, 
        \DATA_OUT_1_48[24]\, \DATA_OUT_1_48[25]\, 
        \DATA_OUT_1_49[0]\, \DATA_OUT_1_49[1]\, 
        \DATA_OUT_1_49[2]\, \DATA_OUT_1_49[3]\, 
        \DATA_OUT_1_49[4]\, \DATA_OUT_1_49[5]\, 
        \DATA_OUT_1_49[6]\, \DATA_OUT_1_49[7]\, 
        \DATA_OUT_1_49[8]\, \DATA_OUT_1_49[9]\, 
        \DATA_OUT_1_49[10]\, \DATA_OUT_1_49[11]\, 
        \DATA_OUT_1_49[12]\, \DATA_OUT_1_49[13]\, 
        \DATA_OUT_1_49[14]\, \DATA_OUT_1_49[15]\, 
        \DATA_OUT_1_49[16]\, \DATA_OUT_1_49[17]\, 
        \DATA_OUT_1_49[18]\, \DATA_OUT_1_49[19]\, 
        \DATA_OUT_1_49[20]\, \DATA_OUT_1_49[21]\, 
        \DATA_OUT_1_49[22]\, \DATA_OUT_1_49[23]\, 
        \DATA_OUT_1_49[24]\, \DATA_OUT_1_49[25]\, 
        \DATA_OUT_1_50[0]\, \DATA_OUT_1_50[1]\, 
        \DATA_OUT_1_50[2]\, \DATA_OUT_1_50[3]\, 
        \DATA_OUT_1_50[4]\, \DATA_OUT_1_50[5]\, 
        \DATA_OUT_1_50[6]\, \DATA_OUT_1_50[7]\, 
        \DATA_OUT_1_50[8]\, \DATA_OUT_1_50[9]\, 
        \DATA_OUT_1_50[10]\, \DATA_OUT_1_50[11]\, 
        \DATA_OUT_1_50[12]\, \DATA_OUT_1_50[13]\, 
        \DATA_OUT_1_50[14]\, \DATA_OUT_1_50[15]\, 
        \DATA_OUT_1_50[16]\, \DATA_OUT_1_50[17]\, 
        \DATA_OUT_1_50[18]\, \DATA_OUT_1_50[19]\, 
        \DATA_OUT_1_50[20]\, \DATA_OUT_1_50[21]\, 
        \DATA_OUT_1_50[22]\, \DATA_OUT_1_50[23]\, 
        \DATA_OUT_1_50[24]\, \DATA_OUT_1_50[25]\, 
        \DATA_OUT_1_51[1]\, \DATA_OUT_1_51[2]\, 
        \DATA_OUT_1_51[3]\, \DATA_OUT_1_51[4]\, 
        \DATA_OUT_1_51[5]\, \DATA_OUT_1_51[6]\, 
        \DATA_OUT_1_51[7]\, \DATA_OUT_1_51[8]\, 
        \DATA_OUT_1_51[9]\, \DATA_OUT_1_51[10]\, 
        \DATA_OUT_1_51[11]\, \DATA_OUT_1_51[12]\, 
        \DATA_OUT_1_51[13]\, \DATA_OUT_1_51[14]\, 
        \DATA_OUT_1_51[15]\, \DATA_OUT_1_51[16]\, 
        \DATA_OUT_1_51[17]\, \DATA_OUT_1_51[18]\, 
        \DATA_OUT_1_51[19]\, \DATA_OUT_1_51[20]\, 
        \DATA_OUT_1_51[21]\, \DATA_OUT_1_51[22]\, 
        \DATA_OUT_1_51[23]\, \DATA_OUT_1_51[24]\, 
        \DATA_OUT_1_51[25]\, \DATA_OR_0_3[0]\, \DATA_OR_0_3[1]\, 
        \DATA_OR_0_3[2]\, \DATA_OR_0_3[3]\, \DATA_OR_0_3[4]\, 
        \DATA_OR_0_3[5]\, \DATA_OR_0_3[6]\, \DATA_OR_0_3[7]\, 
        \DATA_OR_0_3[8]\, \DATA_OR_0_3[9]\, \DATA_OR_0_3[10]\, 
        \DATA_OR_0_3[11]\, \DATA_OR_0_3[12]\, \DATA_OR_0_3[13]\, 
        \DATA_OR_0_3[14]\, \DATA_OR_0_3[15]\, \DATA_OR_0_3[16]\, 
        \DATA_OR_0_3[17]\, \DATA_OR_0_3[18]\, \DATA_OR_0_3[19]\, 
        \DATA_OR_0_3[20]\, \DATA_OR_0_3[21]\, \DATA_OR_0_3[22]\, 
        \DATA_OR_0_3[23]\, \DATA_OR_0_3[24]\, \DATA_OR_0_3[25]\, 
        \DATA_OR_0_0[0]\, \DATA_OR_0_0[1]\, \DATA_OR_0_0[2]\, 
        \DATA_OR_0_0[3]\, \DATA_OR_0_0[4]\, \DATA_OR_0_0[5]\, 
        \DATA_OR_0_0[6]\, \DATA_OR_0_0[7]\, \DATA_OR_0_0[8]\, 
        \DATA_OR_0_0[9]\, \DATA_OR_0_0[10]\, \DATA_OR_0_0[11]\, 
        \DATA_OR_0_0[12]\, \DATA_OR_0_0[13]\, \DATA_OR_0_0[14]\, 
        \DATA_OR_0_0[15]\, \DATA_OR_0_0[16]\, \DATA_OR_0_0[17]\, 
        \DATA_OR_0_0[18]\, \DATA_OR_0_0[19]\, \DATA_OR_0_0[20]\, 
        \DATA_OR_0_0[21]\, \DATA_OR_0_0[22]\, \DATA_OR_0_0[23]\, 
        \DATA_OR_0_0[24]\, \DATA_OR_0_0[25]\, \DATA_OR_0_1[0]\, 
        \DATA_OR_0_1[1]\, \DATA_OR_0_1[2]\, \DATA_OR_0_1[3]\, 
        \DATA_OR_0_1[4]\, \DATA_OR_0_1[5]\, \DATA_OR_0_1[6]\, 
        \DATA_OR_0_1[7]\, \DATA_OR_0_1[8]\, \DATA_OR_0_1[9]\, 
        \DATA_OR_0_1[10]\, \DATA_OR_0_1[11]\, \DATA_OR_0_1[12]\, 
        \DATA_OR_0_1[13]\, \DATA_OR_0_1[14]\, \DATA_OR_0_1[15]\, 
        \DATA_OR_0_1[16]\, \DATA_OR_0_1[17]\, \DATA_OR_0_1[18]\, 
        \DATA_OR_0_1[19]\, \DATA_OR_0_1[20]\, \DATA_OR_0_1[21]\, 
        \DATA_OR_0_1[22]\, \DATA_OR_0_1[23]\, \DATA_OR_0_1[24]\, 
        \DATA_OR_0_1[25]\, \DATA_OR_0_2[0]\, \DATA_OR_0_2[1]\, 
        \DATA_OR_0_2[2]\, \DATA_OR_0_2[3]\, \DATA_OR_0_2[4]\, 
        \DATA_OR_0_2[5]\, \DATA_OR_0_2[6]\, \DATA_OR_0_2[7]\, 
        \DATA_OR_0_2[8]\, \DATA_OR_0_2[9]\, \DATA_OR_0_2[10]\, 
        \DATA_OR_0_2[11]\, \DATA_OR_0_2[12]\, \DATA_OR_0_2[13]\, 
        \DATA_OR_0_2[14]\, \DATA_OR_0_2[15]\, \DATA_OR_0_2[16]\, 
        \DATA_OR_0_2[17]\, \DATA_OR_0_2[18]\, \DATA_OR_0_2[19]\, 
        \DATA_OR_0_2[20]\, \DATA_OR_0_2[21]\, \DATA_OR_0_2[22]\, 
        \DATA_OR_0_2[23]\, \DATA_OR_0_2[24]\, \DATA_OR_0_2[25]\, 
        \DATA_OR_1_0[0]\, \DATA_OR_1_0[1]\, \DATA_OR_1_0[2]\, 
        \DATA_OR_1_0[3]\, \DATA_OR_1_0[4]\, \DATA_OR_1_0[5]\, 
        \DATA_OR_1_0[6]\, \DATA_OR_1_0[7]\, \DATA_OR_1_0[8]\, 
        \DATA_OR_1_0[9]\, \DATA_OR_1_0[10]\, \DATA_OR_1_0[11]\, 
        \DATA_OR_1_0[12]\, \DATA_OR_1_0[13]\, \DATA_OR_1_0[14]\, 
        \DATA_OR_1_0[15]\, \DATA_OR_1_0[16]\, \DATA_OR_1_0[17]\, 
        \DATA_OR_1_0[18]\, \DATA_OR_1_0[19]\, \DATA_OR_1_0[20]\, 
        \DATA_OR_1_0[21]\, \DATA_OR_1_0[22]\, \DATA_OR_1_0[23]\, 
        \DATA_OR_1_0[24]\, \DATA_OR_1_0[25]\, \DATA_OR_1_1[0]\, 
        \DATA_OR_1_1[1]\, \DATA_OR_1_1[2]\, \DATA_OR_1_1[3]\, 
        \DATA_OR_1_1[4]\, \DATA_OR_1_1[5]\, \DATA_OR_1_1[6]\, 
        \DATA_OR_1_1[7]\, \DATA_OR_1_1[8]\, \DATA_OR_1_1[9]\, 
        \DATA_OR_1_1[10]\, \DATA_OR_1_1[11]\, \DATA_OR_1_1[12]\, 
        \DATA_OR_1_1[13]\, \DATA_OR_1_1[14]\, \DATA_OR_1_1[15]\, 
        \DATA_OR_1_1[16]\, \DATA_OR_1_1[17]\, \DATA_OR_1_1[18]\, 
        \DATA_OR_1_1[19]\, \DATA_OR_1_1[20]\, \DATA_OR_1_1[21]\, 
        \DATA_OR_1_1[22]\, \DATA_OR_1_1[23]\, \DATA_OR_1_1[24]\, 
        \DATA_OR_1_1[25]\, \DATA_OR_1_2[0]\, \DATA_OR_1_2[1]\, 
        \DATA_OR_1_2[2]\, \DATA_OR_1_2[3]\, \DATA_OR_1_2[4]\, 
        \DATA_OR_1_2[5]\, \DATA_OR_1_2[6]\, \DATA_OR_1_2[7]\, 
        \DATA_OR_1_2[8]\, \DATA_OR_1_2[9]\, \DATA_OR_1_2[10]\, 
        \DATA_OR_1_2[11]\, \DATA_OR_1_2[12]\, \DATA_OR_1_2[13]\, 
        \DATA_OR_1_2[14]\, \DATA_OR_1_2[15]\, \DATA_OR_1_2[16]\, 
        \DATA_OR_1_2[17]\, \DATA_OR_1_2[18]\, \DATA_OR_1_2[19]\, 
        \DATA_OR_1_2[20]\, \DATA_OR_1_2[21]\, \DATA_OR_1_2[22]\, 
        \DATA_OR_1_2[23]\, \DATA_OR_1_2[24]\, \DATA_OR_1_2[25]\, 
        \DATA_OR_1_3[0]\, \DATA_OR_1_3[1]\, \DATA_OR_1_3[2]\, 
        \DATA_OR_1_3[3]\, \DATA_OR_1_3[4]\, \DATA_OR_1_3[5]\, 
        \DATA_OR_1_3[6]\, \DATA_OR_1_3[7]\, \DATA_OR_1_3[8]\, 
        \DATA_OR_1_3[9]\, \DATA_OR_1_3[10]\, \DATA_OR_1_3[11]\, 
        \DATA_OR_1_3[12]\, \DATA_OR_1_3[13]\, \DATA_OR_1_3[14]\, 
        \DATA_OR_1_3[15]\, \DATA_OR_1_3[16]\, \DATA_OR_1_3[17]\, 
        \DATA_OR_1_3[18]\, \DATA_OR_1_3[19]\, \DATA_OR_1_3[20]\, 
        \DATA_OR_1_3[21]\, \DATA_OR_1_3[22]\, \DATA_OR_1_3[23]\, 
        \DATA_OR_1_3[24]\, \DATA_OR_1_3[25]\, \DATA_OR_1_4[0]\, 
        \DATA_OR_1_4[1]\, \DATA_OR_1_4[2]\, \DATA_OR_1_4[3]\, 
        \DATA_OR_1_4[4]\, \DATA_OR_1_4[5]\, \DATA_OR_1_4[6]\, 
        \DATA_OR_1_4[7]\, \DATA_OR_1_4[8]\, \DATA_OR_1_4[9]\, 
        \DATA_OR_1_4[10]\, \DATA_OR_1_4[11]\, \DATA_OR_1_4[12]\, 
        \DATA_OR_1_4[13]\, \DATA_OR_1_4[14]\, \DATA_OR_1_4[15]\, 
        \DATA_OR_1_4[16]\, \DATA_OR_1_4[17]\, \DATA_OR_1_4[18]\, 
        \DATA_OR_1_4[19]\, \DATA_OR_1_4[20]\, \DATA_OR_1_4[21]\, 
        \DATA_OR_1_4[22]\, \DATA_OR_1_4[23]\, \DATA_OR_1_4[24]\, 
        \DATA_OR_1_4[25]\, \DATA_OR_1_5[0]\, \DATA_OR_1_5[1]\, 
        \DATA_OR_1_5[2]\, \DATA_OR_1_5[3]\, \DATA_OR_1_5[4]\, 
        \DATA_OR_1_5[5]\, \DATA_OR_1_5[6]\, \DATA_OR_1_5[7]\, 
        \DATA_OR_1_5[8]\, \DATA_OR_1_5[9]\, \DATA_OR_1_5[10]\, 
        \DATA_OR_1_5[11]\, \DATA_OR_1_5[12]\, \DATA_OR_1_5[13]\, 
        \DATA_OR_1_5[14]\, \DATA_OR_1_5[15]\, \DATA_OR_1_5[16]\, 
        \DATA_OR_1_5[17]\, \DATA_OR_1_5[18]\, \DATA_OR_1_5[19]\, 
        \DATA_OR_1_5[20]\, \DATA_OR_1_5[21]\, \DATA_OR_1_5[22]\, 
        \DATA_OR_1_5[23]\, \DATA_OR_1_5[24]\, \DATA_OR_1_5[25]\, 
        \DATA_OUT_0_tmp[0]\, \DATA_OUT_0_tmp[1]\, 
        \DATA_OUT_0_tmp[2]\, \DATA_OUT_0_tmp[3]\, 
        \DATA_OUT_0_tmp[4]\, \DATA_OUT_0_tmp[5]\, 
        \DATA_OUT_0_tmp[6]\, \DATA_OUT_0_tmp[7]\, 
        \DATA_OUT_0_tmp[8]\, \DATA_OUT_0_tmp[9]\, 
        \DATA_OUT_0_tmp[10]\, \DATA_OUT_0_tmp[11]\, 
        \DATA_OUT_0_tmp[12]\, \DATA_OUT_0_tmp[13]\, 
        \DATA_OUT_0_tmp[14]\, \DATA_OUT_0_tmp[15]\, 
        \DATA_OUT_0_tmp[16]\, \DATA_OUT_0_tmp[17]\, 
        \DATA_OUT_0_tmp[18]\, \DATA_OUT_0_tmp[19]\, 
        \DATA_OUT_0_tmp[20]\, \DATA_OUT_0_tmp[21]\, 
        \DATA_OUT_0_tmp[22]\, \DATA_OUT_0_tmp[23]\, 
        \DATA_OUT_0_tmp[24]\, \DATA_OUT_0_tmp[25]\, 
        \DATA_OUT_0_tmp[26]\, \DATA_OUT_0_tmp[27]\, 
        \DATA_OUT_0_tmp[28]\, \DATA_OUT_0_tmp[29]\, 
        \DATA_OUT_0_tmp[30]\, \DATA_OUT_0_tmp[31]\, 
        \DATA_OUT_1_tmp[0]\, \DATA_OUT_1_tmp[1]\, 
        \DATA_OUT_1_tmp[2]\, \DATA_OUT_1_tmp[3]\, 
        \DATA_OUT_1_tmp[4]\, \DATA_OUT_1_tmp[5]\, 
        \DATA_OUT_1_tmp[6]\, \DATA_OUT_1_tmp[7]\, 
        \DATA_OUT_1_tmp[8]\, \DATA_OUT_1_tmp[9]\, 
        \DATA_OUT_1_tmp[10]\, \DATA_OUT_1_tmp[11]\, 
        \DATA_OUT_1_tmp[12]\, \DATA_OUT_1_tmp[13]\, 
        \DATA_OUT_1_tmp[14]\, \DATA_OUT_1_tmp[15]\, 
        \DATA_OUT_1_tmp[16]\, \DATA_OUT_1_tmp[17]\, 
        \DATA_OUT_1_tmp[18]\, \DATA_OUT_1_tmp[19]\, 
        \DATA_OUT_1_tmp[20]\, \DATA_OUT_1_tmp[21]\, 
        \DATA_OUT_1_tmp[22]\, \DATA_OUT_1_tmp[23]\, 
        \DATA_OUT_1_tmp[24]\, \DATA_OUT_1_tmp[25]\, 
        \DATA_OUT_1_tmp[26]\, \DATA_OUT_1_tmp[27]\, 
        \DATA_OUT_1_tmp[28]\, \DATA_OUT_1_tmp[29]\, 
        \DATA_OUT_1_tmp[30]\, \DATA_OUT_1_tmp[31]\, 
        \DATA_OUT_2_tmp[1]\, \DATA_OUT_2_tmp[2]\, 
        \DATA_OUT_2_tmp[3]\, \DATA_OUT_2_tmp[4]\, 
        \DATA_OUT_2_tmp[5]\, \DATA_OUT_2_tmp[6]\, 
        \DATA_OUT_2_tmp[7]\, \DATA_OUT_2_tmp[8]\, 
        \DATA_OUT_2_tmp[9]\, \DATA_OUT_2_tmp[10]\, 
        \DATA_OUT_2_tmp[11]\, \DATA_OUT_2_tmp[12]\, 
        \DATA_OUT_2_tmp[13]\, \DATA_OUT_2_tmp[14]\, 
        \DATA_OUT_2_tmp[15]\, \DATA_OUT_2_tmp[16]\, 
        \DATA_OUT_2_tmp[17]\, \DATA_OUT_2_tmp[18]\, 
        \DATA_OUT_2_tmp[19]\, \DATA_OUT_2_tmp[20]\, 
        \DATA_OUT_2_tmp[21]\, \DATA_OUT_2_tmp[22]\, 
        \DATA_OUT_2_tmp[23]\, \DATA_OUT_2_tmp[24]\, 
        \DATA_OUT_2_tmp[25]\, \DATA_OUT_2_tmp[26]\, 
        \DATA_OUT_2_tmp[27]\, \DATA_OUT_2_tmp[28]\, 
        \DATA_OUT_2_tmp[29]\, \DATA_OUT_2_tmp[30]\, 
        \DATA_OUT_2_tmp[31]\, \DATA_OUT_3_tmp[1]\, 
        \DATA_OUT_3_tmp[2]\, \DATA_OUT_3_tmp[3]\, 
        \DATA_OUT_3_tmp[4]\, \DATA_OUT_3_tmp[5]\, 
        \DATA_OUT_3_tmp[6]\, \DATA_OUT_3_tmp[7]\, 
        \DATA_OUT_3_tmp[8]\, \DATA_OUT_3_tmp[9]\, 
        \DATA_OUT_3_tmp[10]\, \DATA_OUT_3_tmp[11]\, 
        \DATA_OUT_3_tmp[12]\, \DATA_OUT_3_tmp[13]\, 
        \DATA_OUT_3_tmp[14]\, \DATA_OUT_3_tmp[15]\, 
        \DATA_OUT_3_tmp[16]\, \DATA_OUT_3_tmp[17]\, 
        \DATA_OUT_3_tmp[18]\, \DATA_OUT_3_tmp[19]\, 
        \DATA_OUT_3_tmp[20]\, \DATA_OUT_3_tmp[21]\, 
        \DATA_OUT_3_tmp[22]\, \DATA_OUT_3_tmp[23]\, 
        \DATA_OUT_3_tmp[24]\, \DATA_OUT_3_tmp[25]\, 
        \DATA_OUT_3_tmp[26]\, \DATA_OUT_3_tmp[27]\, 
        \DATA_OUT_3_tmp[28]\, \DATA_OUT_3_tmp[29]\, 
        \DATA_OUT_3_tmp[30]\, \DATA_OUT_3_tmp[31]\, \VCC\, GND_0, 
        VCC_0 : std_logic;

begin 

    \DATA_IN_1[103]\ <= DATA_IN_1(103);
    TEST_OUT(7) <= \GND\;
    TEST_OUT(6) <= \GND\;
    TEST_OUT(5) <= \GND\;
    TEST_OUT(4) <= \DATA_OUT_2_tmp[0]\;
    TEST_OUT(3) <= \DATA_OUT_3_tmp[0]\;
    TEST_OUT(2) <= \DATA_OUT_1_51[0]\;
    TEST_OUT(1) <= \DATA_OUT_PF_1[103]\;
    TEST_OUT(0) <= \DATA_IN_1[103]\;

    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    Inst_or_array : or_array
      port map(CLK => CLK, RST => RST, DATA_IN_0_0(25) => 
        \DATA_OUT_0_0[25]\, DATA_IN_0_0(24) => \DATA_OUT_0_0[24]\, 
        DATA_IN_0_0(23) => \DATA_OUT_0_0[23]\, DATA_IN_0_0(22)
         => \DATA_OUT_0_0[22]\, DATA_IN_0_0(21) => 
        \DATA_OUT_0_0[21]\, DATA_IN_0_0(20) => \DATA_OUT_0_0[20]\, 
        DATA_IN_0_0(19) => \DATA_OUT_0_0[19]\, DATA_IN_0_0(18)
         => \DATA_OUT_0_0[18]\, DATA_IN_0_0(17) => 
        \DATA_OUT_0_0[17]\, DATA_IN_0_0(16) => \DATA_OUT_0_0[16]\, 
        DATA_IN_0_0(15) => \DATA_OUT_0_0[15]\, DATA_IN_0_0(14)
         => \DATA_OUT_0_0[14]\, DATA_IN_0_0(13) => 
        \DATA_OUT_0_0[13]\, DATA_IN_0_0(12) => \DATA_OUT_0_0[12]\, 
        DATA_IN_0_0(11) => \DATA_OUT_0_0[11]\, DATA_IN_0_0(10)
         => \DATA_OUT_0_0[10]\, DATA_IN_0_0(9) => 
        \DATA_OUT_0_0[9]\, DATA_IN_0_0(8) => \DATA_OUT_0_0[8]\, 
        DATA_IN_0_0(7) => \DATA_OUT_0_0[7]\, DATA_IN_0_0(6) => 
        \DATA_OUT_0_0[6]\, DATA_IN_0_0(5) => \DATA_OUT_0_0[5]\, 
        DATA_IN_0_0(4) => \DATA_OUT_0_0[4]\, DATA_IN_0_0(3) => 
        \DATA_OUT_0_0[3]\, DATA_IN_0_0(2) => \DATA_OUT_0_0[2]\, 
        DATA_IN_0_0(1) => \DATA_OUT_0_0[1]\, DATA_IN_0_0(0) => 
        \DATA_OUT_0_0[0]\, DATA_IN_0_1(25) => \DATA_OUT_0_1[25]\, 
        DATA_IN_0_1(24) => \DATA_OUT_0_1[24]\, DATA_IN_0_1(23)
         => \DATA_OUT_0_1[23]\, DATA_IN_0_1(22) => 
        \DATA_OUT_0_1[22]\, DATA_IN_0_1(21) => \DATA_OUT_0_1[21]\, 
        DATA_IN_0_1(20) => \DATA_OUT_0_1[20]\, DATA_IN_0_1(19)
         => \DATA_OUT_0_1[19]\, DATA_IN_0_1(18) => 
        \DATA_OUT_0_1[18]\, DATA_IN_0_1(17) => \DATA_OUT_0_1[17]\, 
        DATA_IN_0_1(16) => \DATA_OUT_0_1[16]\, DATA_IN_0_1(15)
         => \DATA_OUT_0_1[15]\, DATA_IN_0_1(14) => 
        \DATA_OUT_0_1[14]\, DATA_IN_0_1(13) => \DATA_OUT_0_1[13]\, 
        DATA_IN_0_1(12) => \DATA_OUT_0_1[12]\, DATA_IN_0_1(11)
         => \DATA_OUT_0_1[11]\, DATA_IN_0_1(10) => 
        \DATA_OUT_0_1[10]\, DATA_IN_0_1(9) => \DATA_OUT_0_1[9]\, 
        DATA_IN_0_1(8) => \DATA_OUT_0_1[8]\, DATA_IN_0_1(7) => 
        \DATA_OUT_0_1[7]\, DATA_IN_0_1(6) => \DATA_OUT_0_1[6]\, 
        DATA_IN_0_1(5) => \DATA_OUT_0_1[5]\, DATA_IN_0_1(4) => 
        \DATA_OUT_0_1[4]\, DATA_IN_0_1(3) => \DATA_OUT_0_1[3]\, 
        DATA_IN_0_1(2) => \DATA_OUT_0_1[2]\, DATA_IN_0_1(1) => 
        \DATA_OUT_0_1[1]\, DATA_IN_0_1(0) => \DATA_OUT_0_1[0]\, 
        DATA_IN_0_2(25) => \DATA_OUT_0_2[25]\, DATA_IN_0_2(24)
         => \DATA_OUT_0_2[24]\, DATA_IN_0_2(23) => 
        \DATA_OUT_0_2[23]\, DATA_IN_0_2(22) => \DATA_OUT_0_2[22]\, 
        DATA_IN_0_2(21) => \DATA_OUT_0_2[21]\, DATA_IN_0_2(20)
         => \DATA_OUT_0_2[20]\, DATA_IN_0_2(19) => 
        \DATA_OUT_0_2[19]\, DATA_IN_0_2(18) => \DATA_OUT_0_2[18]\, 
        DATA_IN_0_2(17) => \DATA_OUT_0_2[17]\, DATA_IN_0_2(16)
         => \DATA_OUT_0_2[16]\, DATA_IN_0_2(15) => 
        \DATA_OUT_0_2[15]\, DATA_IN_0_2(14) => \DATA_OUT_0_2[14]\, 
        DATA_IN_0_2(13) => \DATA_OUT_0_2[13]\, DATA_IN_0_2(12)
         => \DATA_OUT_0_2[12]\, DATA_IN_0_2(11) => 
        \DATA_OUT_0_2[11]\, DATA_IN_0_2(10) => \DATA_OUT_0_2[10]\, 
        DATA_IN_0_2(9) => \DATA_OUT_0_2[9]\, DATA_IN_0_2(8) => 
        \DATA_OUT_0_2[8]\, DATA_IN_0_2(7) => \DATA_OUT_0_2[7]\, 
        DATA_IN_0_2(6) => \DATA_OUT_0_2[6]\, DATA_IN_0_2(5) => 
        \DATA_OUT_0_2[5]\, DATA_IN_0_2(4) => \DATA_OUT_0_2[4]\, 
        DATA_IN_0_2(3) => \DATA_OUT_0_2[3]\, DATA_IN_0_2(2) => 
        \DATA_OUT_0_2[2]\, DATA_IN_0_2(1) => \DATA_OUT_0_2[1]\, 
        DATA_IN_0_2(0) => \DATA_OUT_0_2[0]\, DATA_IN_0_3(25) => 
        \DATA_OUT_0_3[25]\, DATA_IN_0_3(24) => \DATA_OUT_0_3[24]\, 
        DATA_IN_0_3(23) => \DATA_OUT_0_3[23]\, DATA_IN_0_3(22)
         => \DATA_OUT_0_3[22]\, DATA_IN_0_3(21) => 
        \DATA_OUT_0_3[21]\, DATA_IN_0_3(20) => \DATA_OUT_0_3[20]\, 
        DATA_IN_0_3(19) => \DATA_OUT_0_3[19]\, DATA_IN_0_3(18)
         => \DATA_OUT_0_3[18]\, DATA_IN_0_3(17) => 
        \DATA_OUT_0_3[17]\, DATA_IN_0_3(16) => \DATA_OUT_0_3[16]\, 
        DATA_IN_0_3(15) => \DATA_OUT_0_3[15]\, DATA_IN_0_3(14)
         => \DATA_OUT_0_3[14]\, DATA_IN_0_3(13) => 
        \DATA_OUT_0_3[13]\, DATA_IN_0_3(12) => \DATA_OUT_0_3[12]\, 
        DATA_IN_0_3(11) => \DATA_OUT_0_3[11]\, DATA_IN_0_3(10)
         => \DATA_OUT_0_3[10]\, DATA_IN_0_3(9) => 
        \DATA_OUT_0_3[9]\, DATA_IN_0_3(8) => \DATA_OUT_0_3[8]\, 
        DATA_IN_0_3(7) => \DATA_OUT_0_3[7]\, DATA_IN_0_3(6) => 
        \DATA_OUT_0_3[6]\, DATA_IN_0_3(5) => \DATA_OUT_0_3[5]\, 
        DATA_IN_0_3(4) => \DATA_OUT_0_3[4]\, DATA_IN_0_3(3) => 
        \DATA_OUT_0_3[3]\, DATA_IN_0_3(2) => \DATA_OUT_0_3[2]\, 
        DATA_IN_0_3(1) => \DATA_OUT_0_3[1]\, DATA_IN_0_3(0) => 
        \DATA_OUT_0_3[0]\, DATA_IN_0_4(25) => \DATA_OUT_0_4[25]\, 
        DATA_IN_0_4(24) => \DATA_OUT_0_4[24]\, DATA_IN_0_4(23)
         => \DATA_OUT_0_4[23]\, DATA_IN_0_4(22) => 
        \DATA_OUT_0_4[22]\, DATA_IN_0_4(21) => \DATA_OUT_0_4[21]\, 
        DATA_IN_0_4(20) => \DATA_OUT_0_4[20]\, DATA_IN_0_4(19)
         => \DATA_OUT_0_4[19]\, DATA_IN_0_4(18) => 
        \DATA_OUT_0_4[18]\, DATA_IN_0_4(17) => \DATA_OUT_0_4[17]\, 
        DATA_IN_0_4(16) => \DATA_OUT_0_4[16]\, DATA_IN_0_4(15)
         => \DATA_OUT_0_4[15]\, DATA_IN_0_4(14) => 
        \DATA_OUT_0_4[14]\, DATA_IN_0_4(13) => \DATA_OUT_0_4[13]\, 
        DATA_IN_0_4(12) => \DATA_OUT_0_4[12]\, DATA_IN_0_4(11)
         => \DATA_OUT_0_4[11]\, DATA_IN_0_4(10) => 
        \DATA_OUT_0_4[10]\, DATA_IN_0_4(9) => \DATA_OUT_0_4[9]\, 
        DATA_IN_0_4(8) => \DATA_OUT_0_4[8]\, DATA_IN_0_4(7) => 
        \DATA_OUT_0_4[7]\, DATA_IN_0_4(6) => \DATA_OUT_0_4[6]\, 
        DATA_IN_0_4(5) => \DATA_OUT_0_4[5]\, DATA_IN_0_4(4) => 
        \DATA_OUT_0_4[4]\, DATA_IN_0_4(3) => \DATA_OUT_0_4[3]\, 
        DATA_IN_0_4(2) => \DATA_OUT_0_4[2]\, DATA_IN_0_4(1) => 
        \DATA_OUT_0_4[1]\, DATA_IN_0_4(0) => \DATA_OUT_0_4[0]\, 
        DATA_IN_0_5(25) => \DATA_OUT_0_5[25]\, DATA_IN_0_5(24)
         => \DATA_OUT_0_5[24]\, DATA_IN_0_5(23) => 
        \DATA_OUT_0_5[23]\, DATA_IN_0_5(22) => \DATA_OUT_0_5[22]\, 
        DATA_IN_0_5(21) => \DATA_OUT_0_5[21]\, DATA_IN_0_5(20)
         => \DATA_OUT_0_5[20]\, DATA_IN_0_5(19) => 
        \DATA_OUT_0_5[19]\, DATA_IN_0_5(18) => \DATA_OUT_0_5[18]\, 
        DATA_IN_0_5(17) => \DATA_OUT_0_5[17]\, DATA_IN_0_5(16)
         => \DATA_OUT_0_5[16]\, DATA_IN_0_5(15) => 
        \DATA_OUT_0_5[15]\, DATA_IN_0_5(14) => \DATA_OUT_0_5[14]\, 
        DATA_IN_0_5(13) => \DATA_OUT_0_5[13]\, DATA_IN_0_5(12)
         => \DATA_OUT_0_5[12]\, DATA_IN_0_5(11) => 
        \DATA_OUT_0_5[11]\, DATA_IN_0_5(10) => \DATA_OUT_0_5[10]\, 
        DATA_IN_0_5(9) => \DATA_OUT_0_5[9]\, DATA_IN_0_5(8) => 
        \DATA_OUT_0_5[8]\, DATA_IN_0_5(7) => \DATA_OUT_0_5[7]\, 
        DATA_IN_0_5(6) => \DATA_OUT_0_5[6]\, DATA_IN_0_5(5) => 
        \DATA_OUT_0_5[5]\, DATA_IN_0_5(4) => \DATA_OUT_0_5[4]\, 
        DATA_IN_0_5(3) => \DATA_OUT_0_5[3]\, DATA_IN_0_5(2) => 
        \DATA_OUT_0_5[2]\, DATA_IN_0_5(1) => \DATA_OUT_0_5[1]\, 
        DATA_IN_0_5(0) => \DATA_OUT_0_5[0]\, DATA_IN_0_6(25) => 
        \DATA_OUT_0_6[25]\, DATA_IN_0_6(24) => \DATA_OUT_0_6[24]\, 
        DATA_IN_0_6(23) => \DATA_OUT_0_6[23]\, DATA_IN_0_6(22)
         => \DATA_OUT_0_6[22]\, DATA_IN_0_6(21) => 
        \DATA_OUT_0_6[21]\, DATA_IN_0_6(20) => \DATA_OUT_0_6[20]\, 
        DATA_IN_0_6(19) => \DATA_OUT_0_6[19]\, DATA_IN_0_6(18)
         => \DATA_OUT_0_6[18]\, DATA_IN_0_6(17) => 
        \DATA_OUT_0_6[17]\, DATA_IN_0_6(16) => \DATA_OUT_0_6[16]\, 
        DATA_IN_0_6(15) => \DATA_OUT_0_6[15]\, DATA_IN_0_6(14)
         => \DATA_OUT_0_6[14]\, DATA_IN_0_6(13) => 
        \DATA_OUT_0_6[13]\, DATA_IN_0_6(12) => \DATA_OUT_0_6[12]\, 
        DATA_IN_0_6(11) => \DATA_OUT_0_6[11]\, DATA_IN_0_6(10)
         => \DATA_OUT_0_6[10]\, DATA_IN_0_6(9) => 
        \DATA_OUT_0_6[9]\, DATA_IN_0_6(8) => \DATA_OUT_0_6[8]\, 
        DATA_IN_0_6(7) => \DATA_OUT_0_6[7]\, DATA_IN_0_6(6) => 
        \DATA_OUT_0_6[6]\, DATA_IN_0_6(5) => \DATA_OUT_0_6[5]\, 
        DATA_IN_0_6(4) => \DATA_OUT_0_6[4]\, DATA_IN_0_6(3) => 
        \DATA_OUT_0_6[3]\, DATA_IN_0_6(2) => \DATA_OUT_0_6[2]\, 
        DATA_IN_0_6(1) => \DATA_OUT_0_6[1]\, DATA_IN_0_6(0) => 
        \DATA_OUT_0_6[0]\, DATA_IN_0_7(25) => \DATA_OUT_0_7[25]\, 
        DATA_IN_0_7(24) => \DATA_OUT_0_7[24]\, DATA_IN_0_7(23)
         => \DATA_OUT_0_7[23]\, DATA_IN_0_7(22) => 
        \DATA_OUT_0_7[22]\, DATA_IN_0_7(21) => \DATA_OUT_0_7[21]\, 
        DATA_IN_0_7(20) => \DATA_OUT_0_7[20]\, DATA_IN_0_7(19)
         => \DATA_OUT_0_7[19]\, DATA_IN_0_7(18) => 
        \DATA_OUT_0_7[18]\, DATA_IN_0_7(17) => \DATA_OUT_0_7[17]\, 
        DATA_IN_0_7(16) => \DATA_OUT_0_7[16]\, DATA_IN_0_7(15)
         => \DATA_OUT_0_7[15]\, DATA_IN_0_7(14) => 
        \DATA_OUT_0_7[14]\, DATA_IN_0_7(13) => \DATA_OUT_0_7[13]\, 
        DATA_IN_0_7(12) => \DATA_OUT_0_7[12]\, DATA_IN_0_7(11)
         => \DATA_OUT_0_7[11]\, DATA_IN_0_7(10) => 
        \DATA_OUT_0_7[10]\, DATA_IN_0_7(9) => \DATA_OUT_0_7[9]\, 
        DATA_IN_0_7(8) => \DATA_OUT_0_7[8]\, DATA_IN_0_7(7) => 
        \DATA_OUT_0_7[7]\, DATA_IN_0_7(6) => \DATA_OUT_0_7[6]\, 
        DATA_IN_0_7(5) => \DATA_OUT_0_7[5]\, DATA_IN_0_7(4) => 
        \DATA_OUT_0_7[4]\, DATA_IN_0_7(3) => \DATA_OUT_0_7[3]\, 
        DATA_IN_0_7(2) => \DATA_OUT_0_7[2]\, DATA_IN_0_7(1) => 
        \DATA_OUT_0_7[1]\, DATA_IN_0_7(0) => \DATA_OUT_0_7[0]\, 
        DATA_IN_0_8(25) => \DATA_OUT_0_8[25]\, DATA_IN_0_8(24)
         => \DATA_OUT_0_8[24]\, DATA_IN_0_8(23) => 
        \DATA_OUT_0_8[23]\, DATA_IN_0_8(22) => \DATA_OUT_0_8[22]\, 
        DATA_IN_0_8(21) => \DATA_OUT_0_8[21]\, DATA_IN_0_8(20)
         => \DATA_OUT_0_8[20]\, DATA_IN_0_8(19) => 
        \DATA_OUT_0_8[19]\, DATA_IN_0_8(18) => \DATA_OUT_0_8[18]\, 
        DATA_IN_0_8(17) => \DATA_OUT_0_8[17]\, DATA_IN_0_8(16)
         => \DATA_OUT_0_8[16]\, DATA_IN_0_8(15) => 
        \DATA_OUT_0_8[15]\, DATA_IN_0_8(14) => \DATA_OUT_0_8[14]\, 
        DATA_IN_0_8(13) => \DATA_OUT_0_8[13]\, DATA_IN_0_8(12)
         => \DATA_OUT_0_8[12]\, DATA_IN_0_8(11) => 
        \DATA_OUT_0_8[11]\, DATA_IN_0_8(10) => \DATA_OUT_0_8[10]\, 
        DATA_IN_0_8(9) => \DATA_OUT_0_8[9]\, DATA_IN_0_8(8) => 
        \DATA_OUT_0_8[8]\, DATA_IN_0_8(7) => \DATA_OUT_0_8[7]\, 
        DATA_IN_0_8(6) => \DATA_OUT_0_8[6]\, DATA_IN_0_8(5) => 
        \DATA_OUT_0_8[5]\, DATA_IN_0_8(4) => \DATA_OUT_0_8[4]\, 
        DATA_IN_0_8(3) => \DATA_OUT_0_8[3]\, DATA_IN_0_8(2) => 
        \DATA_OUT_0_8[2]\, DATA_IN_0_8(1) => \DATA_OUT_0_8[1]\, 
        DATA_IN_0_8(0) => \DATA_OUT_0_8[0]\, DATA_IN_0_9(25) => 
        \DATA_OUT_0_9[25]\, DATA_IN_0_9(24) => \DATA_OUT_0_9[24]\, 
        DATA_IN_0_9(23) => \DATA_OUT_0_9[23]\, DATA_IN_0_9(22)
         => \DATA_OUT_0_9[22]\, DATA_IN_0_9(21) => 
        \DATA_OUT_0_9[21]\, DATA_IN_0_9(20) => \DATA_OUT_0_9[20]\, 
        DATA_IN_0_9(19) => \DATA_OUT_0_9[19]\, DATA_IN_0_9(18)
         => \DATA_OUT_0_9[18]\, DATA_IN_0_9(17) => 
        \DATA_OUT_0_9[17]\, DATA_IN_0_9(16) => \DATA_OUT_0_9[16]\, 
        DATA_IN_0_9(15) => \DATA_OUT_0_9[15]\, DATA_IN_0_9(14)
         => \DATA_OUT_0_9[14]\, DATA_IN_0_9(13) => 
        \DATA_OUT_0_9[13]\, DATA_IN_0_9(12) => \DATA_OUT_0_9[12]\, 
        DATA_IN_0_9(11) => \DATA_OUT_0_9[11]\, DATA_IN_0_9(10)
         => \DATA_OUT_0_9[10]\, DATA_IN_0_9(9) => 
        \DATA_OUT_0_9[9]\, DATA_IN_0_9(8) => \DATA_OUT_0_9[8]\, 
        DATA_IN_0_9(7) => \DATA_OUT_0_9[7]\, DATA_IN_0_9(6) => 
        \DATA_OUT_0_9[6]\, DATA_IN_0_9(5) => \DATA_OUT_0_9[5]\, 
        DATA_IN_0_9(4) => \DATA_OUT_0_9[4]\, DATA_IN_0_9(3) => 
        \DATA_OUT_0_9[3]\, DATA_IN_0_9(2) => \DATA_OUT_0_9[2]\, 
        DATA_IN_0_9(1) => \DATA_OUT_0_9[1]\, DATA_IN_0_9(0) => 
        \DATA_OUT_0_9[0]\, DATA_IN_0_26(25) => 
        \DATA_OUT_0_26[25]\, DATA_IN_0_26(24) => 
        \DATA_OUT_0_26[24]\, DATA_IN_0_26(23) => 
        \DATA_OUT_0_26[23]\, DATA_IN_0_26(22) => 
        \DATA_OUT_0_26[22]\, DATA_IN_0_26(21) => 
        \DATA_OUT_0_26[21]\, DATA_IN_0_26(20) => 
        \DATA_OUT_0_26[20]\, DATA_IN_0_26(19) => 
        \DATA_OUT_0_26[19]\, DATA_IN_0_26(18) => 
        \DATA_OUT_0_26[18]\, DATA_IN_0_26(17) => 
        \DATA_OUT_0_26[17]\, DATA_IN_0_26(16) => 
        \DATA_OUT_0_26[16]\, DATA_IN_0_26(15) => 
        \DATA_OUT_0_26[15]\, DATA_IN_0_26(14) => 
        \DATA_OUT_0_26[14]\, DATA_IN_0_26(13) => 
        \DATA_OUT_0_26[13]\, DATA_IN_0_26(12) => 
        \DATA_OUT_0_26[12]\, DATA_IN_0_26(11) => 
        \DATA_OUT_0_26[11]\, DATA_IN_0_26(10) => 
        \DATA_OUT_0_26[10]\, DATA_IN_0_26(9) => 
        \DATA_OUT_0_26[9]\, DATA_IN_0_26(8) => \DATA_OUT_0_26[8]\, 
        DATA_IN_0_26(7) => \DATA_OUT_0_26[7]\, DATA_IN_0_26(6)
         => \DATA_OUT_0_26[6]\, DATA_IN_0_26(5) => 
        \DATA_OUT_0_26[5]\, DATA_IN_0_26(4) => \DATA_OUT_0_26[4]\, 
        DATA_IN_0_26(3) => \DATA_OUT_0_26[3]\, DATA_IN_0_26(2)
         => \DATA_OUT_0_26[2]\, DATA_IN_0_26(1) => 
        \DATA_OUT_0_26[1]\, DATA_IN_0_26(0) => \DATA_OUT_0_26[0]\, 
        DATA_IN_0_27(25) => \DATA_OUT_0_27[25]\, DATA_IN_0_27(24)
         => \DATA_OUT_0_27[24]\, DATA_IN_0_27(23) => 
        \DATA_OUT_0_27[23]\, DATA_IN_0_27(22) => 
        \DATA_OUT_0_27[22]\, DATA_IN_0_27(21) => 
        \DATA_OUT_0_27[21]\, DATA_IN_0_27(20) => 
        \DATA_OUT_0_27[20]\, DATA_IN_0_27(19) => 
        \DATA_OUT_0_27[19]\, DATA_IN_0_27(18) => 
        \DATA_OUT_0_27[18]\, DATA_IN_0_27(17) => 
        \DATA_OUT_0_27[17]\, DATA_IN_0_27(16) => 
        \DATA_OUT_0_27[16]\, DATA_IN_0_27(15) => 
        \DATA_OUT_0_27[15]\, DATA_IN_0_27(14) => 
        \DATA_OUT_0_27[14]\, DATA_IN_0_27(13) => 
        \DATA_OUT_0_27[13]\, DATA_IN_0_27(12) => 
        \DATA_OUT_0_27[12]\, DATA_IN_0_27(11) => 
        \DATA_OUT_0_27[11]\, DATA_IN_0_27(10) => 
        \DATA_OUT_0_27[10]\, DATA_IN_0_27(9) => 
        \DATA_OUT_0_27[9]\, DATA_IN_0_27(8) => \DATA_OUT_0_27[8]\, 
        DATA_IN_0_27(7) => \DATA_OUT_0_27[7]\, DATA_IN_0_27(6)
         => \DATA_OUT_0_27[6]\, DATA_IN_0_27(5) => 
        \DATA_OUT_0_27[5]\, DATA_IN_0_27(4) => \DATA_OUT_0_27[4]\, 
        DATA_IN_0_27(3) => \DATA_OUT_0_27[3]\, DATA_IN_0_27(2)
         => \DATA_OUT_0_27[2]\, DATA_IN_0_27(1) => 
        \DATA_OUT_0_27[1]\, DATA_IN_0_27(0) => \DATA_OUT_0_27[0]\, 
        DATA_IN_0_28(25) => \DATA_OUT_0_28[25]\, DATA_IN_0_28(24)
         => \DATA_OUT_0_28[24]\, DATA_IN_0_28(23) => 
        \DATA_OUT_0_28[23]\, DATA_IN_0_28(22) => 
        \DATA_OUT_0_28[22]\, DATA_IN_0_28(21) => 
        \DATA_OUT_0_28[21]\, DATA_IN_0_28(20) => 
        \DATA_OUT_0_28[20]\, DATA_IN_0_28(19) => 
        \DATA_OUT_0_28[19]\, DATA_IN_0_28(18) => 
        \DATA_OUT_0_28[18]\, DATA_IN_0_28(17) => 
        \DATA_OUT_0_28[17]\, DATA_IN_0_28(16) => 
        \DATA_OUT_0_28[16]\, DATA_IN_0_28(15) => 
        \DATA_OUT_0_28[15]\, DATA_IN_0_28(14) => 
        \DATA_OUT_0_28[14]\, DATA_IN_0_28(13) => 
        \DATA_OUT_0_28[13]\, DATA_IN_0_28(12) => 
        \DATA_OUT_0_28[12]\, DATA_IN_0_28(11) => 
        \DATA_OUT_0_28[11]\, DATA_IN_0_28(10) => 
        \DATA_OUT_0_28[10]\, DATA_IN_0_28(9) => 
        \DATA_OUT_0_28[9]\, DATA_IN_0_28(8) => \DATA_OUT_0_28[8]\, 
        DATA_IN_0_28(7) => \DATA_OUT_0_28[7]\, DATA_IN_0_28(6)
         => \DATA_OUT_0_28[6]\, DATA_IN_0_28(5) => 
        \DATA_OUT_0_28[5]\, DATA_IN_0_28(4) => \DATA_OUT_0_28[4]\, 
        DATA_IN_0_28(3) => \DATA_OUT_0_28[3]\, DATA_IN_0_28(2)
         => \DATA_OUT_0_28[2]\, DATA_IN_0_28(1) => 
        \DATA_OUT_0_28[1]\, DATA_IN_0_28(0) => \DATA_OUT_0_28[0]\, 
        DATA_IN_0_29(25) => \DATA_OUT_0_29[25]\, DATA_IN_0_29(24)
         => \DATA_OUT_0_29[24]\, DATA_IN_0_29(23) => 
        \DATA_OUT_0_29[23]\, DATA_IN_0_29(22) => 
        \DATA_OUT_0_29[22]\, DATA_IN_0_29(21) => 
        \DATA_OUT_0_29[21]\, DATA_IN_0_29(20) => 
        \DATA_OUT_0_29[20]\, DATA_IN_0_29(19) => 
        \DATA_OUT_0_29[19]\, DATA_IN_0_29(18) => 
        \DATA_OUT_0_29[18]\, DATA_IN_0_29(17) => 
        \DATA_OUT_0_29[17]\, DATA_IN_0_29(16) => 
        \DATA_OUT_0_29[16]\, DATA_IN_0_29(15) => 
        \DATA_OUT_0_29[15]\, DATA_IN_0_29(14) => 
        \DATA_OUT_0_29[14]\, DATA_IN_0_29(13) => 
        \DATA_OUT_0_29[13]\, DATA_IN_0_29(12) => 
        \DATA_OUT_0_29[12]\, DATA_IN_0_29(11) => 
        \DATA_OUT_0_29[11]\, DATA_IN_0_29(10) => 
        \DATA_OUT_0_29[10]\, DATA_IN_0_29(9) => 
        \DATA_OUT_0_29[9]\, DATA_IN_0_29(8) => \DATA_OUT_0_29[8]\, 
        DATA_IN_0_29(7) => \DATA_OUT_0_29[7]\, DATA_IN_0_29(6)
         => \DATA_OUT_0_29[6]\, DATA_IN_0_29(5) => 
        \DATA_OUT_0_29[5]\, DATA_IN_0_29(4) => \DATA_OUT_0_29[4]\, 
        DATA_IN_0_29(3) => \DATA_OUT_0_29[3]\, DATA_IN_0_29(2)
         => \DATA_OUT_0_29[2]\, DATA_IN_0_29(1) => 
        \DATA_OUT_0_29[1]\, DATA_IN_0_29(0) => \DATA_OUT_0_29[0]\, 
        DATA_IN_0_30(25) => \DATA_OUT_0_30[25]\, DATA_IN_0_30(24)
         => \DATA_OUT_0_30[24]\, DATA_IN_0_30(23) => 
        \DATA_OUT_0_30[23]\, DATA_IN_0_30(22) => 
        \DATA_OUT_0_30[22]\, DATA_IN_0_30(21) => 
        \DATA_OUT_0_30[21]\, DATA_IN_0_30(20) => 
        \DATA_OUT_0_30[20]\, DATA_IN_0_30(19) => 
        \DATA_OUT_0_30[19]\, DATA_IN_0_30(18) => 
        \DATA_OUT_0_30[18]\, DATA_IN_0_30(17) => 
        \DATA_OUT_0_30[17]\, DATA_IN_0_30(16) => 
        \DATA_OUT_0_30[16]\, DATA_IN_0_30(15) => 
        \DATA_OUT_0_30[15]\, DATA_IN_0_30(14) => 
        \DATA_OUT_0_30[14]\, DATA_IN_0_30(13) => 
        \DATA_OUT_0_30[13]\, DATA_IN_0_30(12) => 
        \DATA_OUT_0_30[12]\, DATA_IN_0_30(11) => 
        \DATA_OUT_0_30[11]\, DATA_IN_0_30(10) => 
        \DATA_OUT_0_30[10]\, DATA_IN_0_30(9) => 
        \DATA_OUT_0_30[9]\, DATA_IN_0_30(8) => \DATA_OUT_0_30[8]\, 
        DATA_IN_0_30(7) => \DATA_OUT_0_30[7]\, DATA_IN_0_30(6)
         => \DATA_OUT_0_30[6]\, DATA_IN_0_30(5) => 
        \DATA_OUT_0_30[5]\, DATA_IN_0_30(4) => \DATA_OUT_0_30[4]\, 
        DATA_IN_0_30(3) => \DATA_OUT_0_30[3]\, DATA_IN_0_30(2)
         => \DATA_OUT_0_30[2]\, DATA_IN_0_30(1) => 
        \DATA_OUT_0_30[1]\, DATA_IN_0_30(0) => \DATA_OUT_0_30[0]\, 
        DATA_IN_0_31(25) => \DATA_OUT_0_31[25]\, DATA_IN_0_31(24)
         => \DATA_OUT_0_31[24]\, DATA_IN_0_31(23) => 
        \DATA_OUT_0_31[23]\, DATA_IN_0_31(22) => 
        \DATA_OUT_0_31[22]\, DATA_IN_0_31(21) => 
        \DATA_OUT_0_31[21]\, DATA_IN_0_31(20) => 
        \DATA_OUT_0_31[20]\, DATA_IN_0_31(19) => 
        \DATA_OUT_0_31[19]\, DATA_IN_0_31(18) => 
        \DATA_OUT_0_31[18]\, DATA_IN_0_31(17) => 
        \DATA_OUT_0_31[17]\, DATA_IN_0_31(16) => 
        \DATA_OUT_0_31[16]\, DATA_IN_0_31(15) => 
        \DATA_OUT_0_31[15]\, DATA_IN_0_31(14) => 
        \DATA_OUT_0_31[14]\, DATA_IN_0_31(13) => 
        \DATA_OUT_0_31[13]\, DATA_IN_0_31(12) => 
        \DATA_OUT_0_31[12]\, DATA_IN_0_31(11) => 
        \DATA_OUT_0_31[11]\, DATA_IN_0_31(10) => 
        \DATA_OUT_0_31[10]\, DATA_IN_0_31(9) => 
        \DATA_OUT_0_31[9]\, DATA_IN_0_31(8) => \DATA_OUT_0_31[8]\, 
        DATA_IN_0_31(7) => \DATA_OUT_0_31[7]\, DATA_IN_0_31(6)
         => \DATA_OUT_0_31[6]\, DATA_IN_0_31(5) => 
        \DATA_OUT_0_31[5]\, DATA_IN_0_31(4) => \DATA_OUT_0_31[4]\, 
        DATA_IN_0_31(3) => \DATA_OUT_0_31[3]\, DATA_IN_0_31(2)
         => \DATA_OUT_0_31[2]\, DATA_IN_0_31(1) => 
        \DATA_OUT_0_31[1]\, DATA_IN_0_31(0) => \DATA_OUT_0_31[0]\, 
        DATA_IN_0_32(25) => \DATA_OUT_0_32[25]\, DATA_IN_0_32(24)
         => \DATA_OUT_0_32[24]\, DATA_IN_0_32(23) => 
        \DATA_OUT_0_32[23]\, DATA_IN_0_32(22) => 
        \DATA_OUT_0_32[22]\, DATA_IN_0_32(21) => 
        \DATA_OUT_0_32[21]\, DATA_IN_0_32(20) => 
        \DATA_OUT_0_32[20]\, DATA_IN_0_32(19) => 
        \DATA_OUT_0_32[19]\, DATA_IN_0_32(18) => 
        \DATA_OUT_0_32[18]\, DATA_IN_0_32(17) => 
        \DATA_OUT_0_32[17]\, DATA_IN_0_32(16) => 
        \DATA_OUT_0_32[16]\, DATA_IN_0_32(15) => 
        \DATA_OUT_0_32[15]\, DATA_IN_0_32(14) => 
        \DATA_OUT_0_32[14]\, DATA_IN_0_32(13) => 
        \DATA_OUT_0_32[13]\, DATA_IN_0_32(12) => 
        \DATA_OUT_0_32[12]\, DATA_IN_0_32(11) => 
        \DATA_OUT_0_32[11]\, DATA_IN_0_32(10) => 
        \DATA_OUT_0_32[10]\, DATA_IN_0_32(9) => 
        \DATA_OUT_0_32[9]\, DATA_IN_0_32(8) => \DATA_OUT_0_32[8]\, 
        DATA_IN_0_32(7) => \DATA_OUT_0_32[7]\, DATA_IN_0_32(6)
         => \DATA_OUT_0_32[6]\, DATA_IN_0_32(5) => 
        \DATA_OUT_0_32[5]\, DATA_IN_0_32(4) => \DATA_OUT_0_32[4]\, 
        DATA_IN_0_32(3) => \DATA_OUT_0_32[3]\, DATA_IN_0_32(2)
         => \DATA_OUT_0_32[2]\, DATA_IN_0_32(1) => 
        \DATA_OUT_0_32[1]\, DATA_IN_0_32(0) => \DATA_OUT_0_32[0]\, 
        DATA_IN_0_33(25) => \DATA_OUT_0_33[25]\, DATA_IN_0_33(24)
         => \DATA_OUT_0_33[24]\, DATA_IN_0_33(23) => 
        \DATA_OUT_0_33[23]\, DATA_IN_0_33(22) => 
        \DATA_OUT_0_33[22]\, DATA_IN_0_33(21) => 
        \DATA_OUT_0_33[21]\, DATA_IN_0_33(20) => 
        \DATA_OUT_0_33[20]\, DATA_IN_0_33(19) => 
        \DATA_OUT_0_33[19]\, DATA_IN_0_33(18) => 
        \DATA_OUT_0_33[18]\, DATA_IN_0_33(17) => 
        \DATA_OUT_0_33[17]\, DATA_IN_0_33(16) => 
        \DATA_OUT_0_33[16]\, DATA_IN_0_33(15) => 
        \DATA_OUT_0_33[15]\, DATA_IN_0_33(14) => 
        \DATA_OUT_0_33[14]\, DATA_IN_0_33(13) => 
        \DATA_OUT_0_33[13]\, DATA_IN_0_33(12) => 
        \DATA_OUT_0_33[12]\, DATA_IN_0_33(11) => 
        \DATA_OUT_0_33[11]\, DATA_IN_0_33(10) => 
        \DATA_OUT_0_33[10]\, DATA_IN_0_33(9) => 
        \DATA_OUT_0_33[9]\, DATA_IN_0_33(8) => \DATA_OUT_0_33[8]\, 
        DATA_IN_0_33(7) => \DATA_OUT_0_33[7]\, DATA_IN_0_33(6)
         => \DATA_OUT_0_33[6]\, DATA_IN_0_33(5) => 
        \DATA_OUT_0_33[5]\, DATA_IN_0_33(4) => \DATA_OUT_0_33[4]\, 
        DATA_IN_0_33(3) => \DATA_OUT_0_33[3]\, DATA_IN_0_33(2)
         => \DATA_OUT_0_33[2]\, DATA_IN_0_33(1) => 
        \DATA_OUT_0_33[1]\, DATA_IN_0_33(0) => \DATA_OUT_0_33[0]\, 
        DATA_IN_0_34(25) => \DATA_OUT_0_34[25]\, DATA_IN_0_34(24)
         => \DATA_OUT_0_34[24]\, DATA_IN_0_34(23) => 
        \DATA_OUT_0_34[23]\, DATA_IN_0_34(22) => 
        \DATA_OUT_0_34[22]\, DATA_IN_0_34(21) => 
        \DATA_OUT_0_34[21]\, DATA_IN_0_34(20) => 
        \DATA_OUT_0_34[20]\, DATA_IN_0_34(19) => 
        \DATA_OUT_0_34[19]\, DATA_IN_0_34(18) => 
        \DATA_OUT_0_34[18]\, DATA_IN_0_34(17) => 
        \DATA_OUT_0_34[17]\, DATA_IN_0_34(16) => 
        \DATA_OUT_0_34[16]\, DATA_IN_0_34(15) => 
        \DATA_OUT_0_34[15]\, DATA_IN_0_34(14) => 
        \DATA_OUT_0_34[14]\, DATA_IN_0_34(13) => 
        \DATA_OUT_0_34[13]\, DATA_IN_0_34(12) => 
        \DATA_OUT_0_34[12]\, DATA_IN_0_34(11) => 
        \DATA_OUT_0_34[11]\, DATA_IN_0_34(10) => 
        \DATA_OUT_0_34[10]\, DATA_IN_0_34(9) => 
        \DATA_OUT_0_34[9]\, DATA_IN_0_34(8) => \DATA_OUT_0_34[8]\, 
        DATA_IN_0_34(7) => \DATA_OUT_0_34[7]\, DATA_IN_0_34(6)
         => \DATA_OUT_0_34[6]\, DATA_IN_0_34(5) => 
        \DATA_OUT_0_34[5]\, DATA_IN_0_34(4) => \DATA_OUT_0_34[4]\, 
        DATA_IN_0_34(3) => \DATA_OUT_0_34[3]\, DATA_IN_0_34(2)
         => \DATA_OUT_0_34[2]\, DATA_IN_0_34(1) => 
        \DATA_OUT_0_34[1]\, DATA_IN_0_34(0) => \DATA_OUT_0_34[0]\, 
        DATA_IN_0_35(25) => \DATA_OUT_0_35[25]\, DATA_IN_0_35(24)
         => \DATA_OUT_0_35[24]\, DATA_IN_0_35(23) => 
        \DATA_OUT_0_35[23]\, DATA_IN_0_35(22) => 
        \DATA_OUT_0_35[22]\, DATA_IN_0_35(21) => 
        \DATA_OUT_0_35[21]\, DATA_IN_0_35(20) => 
        \DATA_OUT_0_35[20]\, DATA_IN_0_35(19) => 
        \DATA_OUT_0_35[19]\, DATA_IN_0_35(18) => 
        \DATA_OUT_0_35[18]\, DATA_IN_0_35(17) => 
        \DATA_OUT_0_35[17]\, DATA_IN_0_35(16) => 
        \DATA_OUT_0_35[16]\, DATA_IN_0_35(15) => 
        \DATA_OUT_0_35[15]\, DATA_IN_0_35(14) => 
        \DATA_OUT_0_35[14]\, DATA_IN_0_35(13) => 
        \DATA_OUT_0_35[13]\, DATA_IN_0_35(12) => 
        \DATA_OUT_0_35[12]\, DATA_IN_0_35(11) => 
        \DATA_OUT_0_35[11]\, DATA_IN_0_35(10) => 
        \DATA_OUT_0_35[10]\, DATA_IN_0_35(9) => 
        \DATA_OUT_0_35[9]\, DATA_IN_0_35(8) => \DATA_OUT_0_35[8]\, 
        DATA_IN_0_35(7) => \DATA_OUT_0_35[7]\, DATA_IN_0_35(6)
         => \DATA_OUT_0_35[6]\, DATA_IN_0_35(5) => 
        \DATA_OUT_0_35[5]\, DATA_IN_0_35(4) => \DATA_OUT_0_35[4]\, 
        DATA_IN_0_35(3) => \DATA_OUT_0_35[3]\, DATA_IN_0_35(2)
         => \DATA_OUT_0_35[2]\, DATA_IN_0_35(1) => 
        \DATA_OUT_0_35[1]\, DATA_IN_0_35(0) => \DATA_OUT_0_35[0]\, 
        DATA_IN_0_36(25) => \DATA_OUT_0_36[25]\, DATA_IN_0_36(24)
         => \DATA_OUT_0_36[24]\, DATA_IN_0_36(23) => 
        \DATA_OUT_0_36[23]\, DATA_IN_0_36(22) => 
        \DATA_OUT_0_36[22]\, DATA_IN_0_36(21) => 
        \DATA_OUT_0_36[21]\, DATA_IN_0_36(20) => 
        \DATA_OUT_0_36[20]\, DATA_IN_0_36(19) => 
        \DATA_OUT_0_36[19]\, DATA_IN_0_36(18) => 
        \DATA_OUT_0_36[18]\, DATA_IN_0_36(17) => 
        \DATA_OUT_0_36[17]\, DATA_IN_0_36(16) => 
        \DATA_OUT_0_36[16]\, DATA_IN_0_36(15) => 
        \DATA_OUT_0_36[15]\, DATA_IN_0_36(14) => 
        \DATA_OUT_0_36[14]\, DATA_IN_0_36(13) => 
        \DATA_OUT_0_36[13]\, DATA_IN_0_36(12) => 
        \DATA_OUT_0_36[12]\, DATA_IN_0_36(11) => 
        \DATA_OUT_0_36[11]\, DATA_IN_0_36(10) => 
        \DATA_OUT_0_36[10]\, DATA_IN_0_36(9) => 
        \DATA_OUT_0_36[9]\, DATA_IN_0_36(8) => \DATA_OUT_0_36[8]\, 
        DATA_IN_0_36(7) => \DATA_OUT_0_36[7]\, DATA_IN_0_36(6)
         => \DATA_OUT_0_36[6]\, DATA_IN_0_36(5) => 
        \DATA_OUT_0_36[5]\, DATA_IN_0_36(4) => \DATA_OUT_0_36[4]\, 
        DATA_IN_0_36(3) => \DATA_OUT_0_36[3]\, DATA_IN_0_36(2)
         => \DATA_OUT_0_36[2]\, DATA_IN_0_36(1) => 
        \DATA_OUT_0_36[1]\, DATA_IN_0_36(0) => \DATA_OUT_0_36[0]\, 
        DATA_IN_0_37(25) => \DATA_OUT_0_37[25]\, DATA_IN_0_37(24)
         => \DATA_OUT_0_37[24]\, DATA_IN_0_37(23) => 
        \DATA_OUT_0_37[23]\, DATA_IN_0_37(22) => 
        \DATA_OUT_0_37[22]\, DATA_IN_0_37(21) => 
        \DATA_OUT_0_37[21]\, DATA_IN_0_37(20) => 
        \DATA_OUT_0_37[20]\, DATA_IN_0_37(19) => 
        \DATA_OUT_0_37[19]\, DATA_IN_0_37(18) => 
        \DATA_OUT_0_37[18]\, DATA_IN_0_37(17) => 
        \DATA_OUT_0_37[17]\, DATA_IN_0_37(16) => 
        \DATA_OUT_0_37[16]\, DATA_IN_0_37(15) => 
        \DATA_OUT_0_37[15]\, DATA_IN_0_37(14) => 
        \DATA_OUT_0_37[14]\, DATA_IN_0_37(13) => 
        \DATA_OUT_0_37[13]\, DATA_IN_0_37(12) => 
        \DATA_OUT_0_37[12]\, DATA_IN_0_37(11) => 
        \DATA_OUT_0_37[11]\, DATA_IN_0_37(10) => 
        \DATA_OUT_0_37[10]\, DATA_IN_0_37(9) => 
        \DATA_OUT_0_37[9]\, DATA_IN_0_37(8) => \DATA_OUT_0_37[8]\, 
        DATA_IN_0_37(7) => \DATA_OUT_0_37[7]\, DATA_IN_0_37(6)
         => \DATA_OUT_0_37[6]\, DATA_IN_0_37(5) => 
        \DATA_OUT_0_37[5]\, DATA_IN_0_37(4) => \DATA_OUT_0_37[4]\, 
        DATA_IN_0_37(3) => \DATA_OUT_0_37[3]\, DATA_IN_0_37(2)
         => \DATA_OUT_0_37[2]\, DATA_IN_0_37(1) => 
        \DATA_OUT_0_37[1]\, DATA_IN_0_37(0) => \DATA_OUT_0_37[0]\, 
        DATA_IN_0_38(25) => \DATA_OUT_0_38[25]\, DATA_IN_0_38(24)
         => \DATA_OUT_0_38[24]\, DATA_IN_0_38(23) => 
        \DATA_OUT_0_38[23]\, DATA_IN_0_38(22) => 
        \DATA_OUT_0_38[22]\, DATA_IN_0_38(21) => 
        \DATA_OUT_0_38[21]\, DATA_IN_0_38(20) => 
        \DATA_OUT_0_38[20]\, DATA_IN_0_38(19) => 
        \DATA_OUT_0_38[19]\, DATA_IN_0_38(18) => 
        \DATA_OUT_0_38[18]\, DATA_IN_0_38(17) => 
        \DATA_OUT_0_38[17]\, DATA_IN_0_38(16) => 
        \DATA_OUT_0_38[16]\, DATA_IN_0_38(15) => 
        \DATA_OUT_0_38[15]\, DATA_IN_0_38(14) => 
        \DATA_OUT_0_38[14]\, DATA_IN_0_38(13) => 
        \DATA_OUT_0_38[13]\, DATA_IN_0_38(12) => 
        \DATA_OUT_0_38[12]\, DATA_IN_0_38(11) => 
        \DATA_OUT_0_38[11]\, DATA_IN_0_38(10) => 
        \DATA_OUT_0_38[10]\, DATA_IN_0_38(9) => 
        \DATA_OUT_0_38[9]\, DATA_IN_0_38(8) => \DATA_OUT_0_38[8]\, 
        DATA_IN_0_38(7) => \DATA_OUT_0_38[7]\, DATA_IN_0_38(6)
         => \DATA_OUT_0_38[6]\, DATA_IN_0_38(5) => 
        \DATA_OUT_0_38[5]\, DATA_IN_0_38(4) => \DATA_OUT_0_38[4]\, 
        DATA_IN_0_38(3) => \DATA_OUT_0_38[3]\, DATA_IN_0_38(2)
         => \DATA_OUT_0_38[2]\, DATA_IN_0_38(1) => 
        \DATA_OUT_0_38[1]\, DATA_IN_0_38(0) => \DATA_OUT_0_38[0]\, 
        DATA_IN_0_39(25) => \DATA_OUT_0_39[25]\, DATA_IN_0_39(24)
         => \DATA_OUT_0_39[24]\, DATA_IN_0_39(23) => 
        \DATA_OUT_0_39[23]\, DATA_IN_0_39(22) => 
        \DATA_OUT_0_39[22]\, DATA_IN_0_39(21) => 
        \DATA_OUT_0_39[21]\, DATA_IN_0_39(20) => 
        \DATA_OUT_0_39[20]\, DATA_IN_0_39(19) => 
        \DATA_OUT_0_39[19]\, DATA_IN_0_39(18) => 
        \DATA_OUT_0_39[18]\, DATA_IN_0_39(17) => 
        \DATA_OUT_0_39[17]\, DATA_IN_0_39(16) => 
        \DATA_OUT_0_39[16]\, DATA_IN_0_39(15) => 
        \DATA_OUT_0_39[15]\, DATA_IN_0_39(14) => 
        \DATA_OUT_0_39[14]\, DATA_IN_0_39(13) => 
        \DATA_OUT_0_39[13]\, DATA_IN_0_39(12) => 
        \DATA_OUT_0_39[12]\, DATA_IN_0_39(11) => 
        \DATA_OUT_0_39[11]\, DATA_IN_0_39(10) => 
        \DATA_OUT_0_39[10]\, DATA_IN_0_39(9) => 
        \DATA_OUT_0_39[9]\, DATA_IN_0_39(8) => \DATA_OUT_0_39[8]\, 
        DATA_IN_0_39(7) => \DATA_OUT_0_39[7]\, DATA_IN_0_39(6)
         => \DATA_OUT_0_39[6]\, DATA_IN_0_39(5) => 
        \DATA_OUT_0_39[5]\, DATA_IN_0_39(4) => \DATA_OUT_0_39[4]\, 
        DATA_IN_0_39(3) => \DATA_OUT_0_39[3]\, DATA_IN_0_39(2)
         => \DATA_OUT_0_39[2]\, DATA_IN_0_39(1) => 
        \DATA_OUT_0_39[1]\, DATA_IN_0_39(0) => \DATA_OUT_0_39[0]\, 
        DATA_IN_0_40(25) => \DATA_OUT_0_40[25]\, DATA_IN_0_40(24)
         => \DATA_OUT_0_40[24]\, DATA_IN_0_40(23) => 
        \DATA_OUT_0_40[23]\, DATA_IN_0_40(22) => 
        \DATA_OUT_0_40[22]\, DATA_IN_0_40(21) => 
        \DATA_OUT_0_40[21]\, DATA_IN_0_40(20) => 
        \DATA_OUT_0_40[20]\, DATA_IN_0_40(19) => 
        \DATA_OUT_0_40[19]\, DATA_IN_0_40(18) => 
        \DATA_OUT_0_40[18]\, DATA_IN_0_40(17) => 
        \DATA_OUT_0_40[17]\, DATA_IN_0_40(16) => 
        \DATA_OUT_0_40[16]\, DATA_IN_0_40(15) => 
        \DATA_OUT_0_40[15]\, DATA_IN_0_40(14) => 
        \DATA_OUT_0_40[14]\, DATA_IN_0_40(13) => 
        \DATA_OUT_0_40[13]\, DATA_IN_0_40(12) => 
        \DATA_OUT_0_40[12]\, DATA_IN_0_40(11) => 
        \DATA_OUT_0_40[11]\, DATA_IN_0_40(10) => 
        \DATA_OUT_0_40[10]\, DATA_IN_0_40(9) => 
        \DATA_OUT_0_40[9]\, DATA_IN_0_40(8) => \DATA_OUT_0_40[8]\, 
        DATA_IN_0_40(7) => \DATA_OUT_0_40[7]\, DATA_IN_0_40(6)
         => \DATA_OUT_0_40[6]\, DATA_IN_0_40(5) => 
        \DATA_OUT_0_40[5]\, DATA_IN_0_40(4) => \DATA_OUT_0_40[4]\, 
        DATA_IN_0_40(3) => \DATA_OUT_0_40[3]\, DATA_IN_0_40(2)
         => \DATA_OUT_0_40[2]\, DATA_IN_0_40(1) => 
        \DATA_OUT_0_40[1]\, DATA_IN_0_40(0) => \DATA_OUT_0_40[0]\, 
        DATA_IN_0_41(25) => \DATA_OUT_0_41[25]\, DATA_IN_0_41(24)
         => \DATA_OUT_0_41[24]\, DATA_IN_0_41(23) => 
        \DATA_OUT_0_41[23]\, DATA_IN_0_41(22) => 
        \DATA_OUT_0_41[22]\, DATA_IN_0_41(21) => 
        \DATA_OUT_0_41[21]\, DATA_IN_0_41(20) => 
        \DATA_OUT_0_41[20]\, DATA_IN_0_41(19) => 
        \DATA_OUT_0_41[19]\, DATA_IN_0_41(18) => 
        \DATA_OUT_0_41[18]\, DATA_IN_0_41(17) => 
        \DATA_OUT_0_41[17]\, DATA_IN_0_41(16) => 
        \DATA_OUT_0_41[16]\, DATA_IN_0_41(15) => 
        \DATA_OUT_0_41[15]\, DATA_IN_0_41(14) => 
        \DATA_OUT_0_41[14]\, DATA_IN_0_41(13) => 
        \DATA_OUT_0_41[13]\, DATA_IN_0_41(12) => 
        \DATA_OUT_0_41[12]\, DATA_IN_0_41(11) => 
        \DATA_OUT_0_41[11]\, DATA_IN_0_41(10) => 
        \DATA_OUT_0_41[10]\, DATA_IN_0_41(9) => 
        \DATA_OUT_0_41[9]\, DATA_IN_0_41(8) => \DATA_OUT_0_41[8]\, 
        DATA_IN_0_41(7) => \DATA_OUT_0_41[7]\, DATA_IN_0_41(6)
         => \DATA_OUT_0_41[6]\, DATA_IN_0_41(5) => 
        \DATA_OUT_0_41[5]\, DATA_IN_0_41(4) => \DATA_OUT_0_41[4]\, 
        DATA_IN_0_41(3) => \DATA_OUT_0_41[3]\, DATA_IN_0_41(2)
         => \DATA_OUT_0_41[2]\, DATA_IN_0_41(1) => 
        \DATA_OUT_0_41[1]\, DATA_IN_0_41(0) => \DATA_OUT_0_41[0]\, 
        DATA_IN_0_42(25) => \DATA_OUT_0_42[25]\, DATA_IN_0_42(24)
         => \DATA_OUT_0_42[24]\, DATA_IN_0_42(23) => 
        \DATA_OUT_0_42[23]\, DATA_IN_0_42(22) => 
        \DATA_OUT_0_42[22]\, DATA_IN_0_42(21) => 
        \DATA_OUT_0_42[21]\, DATA_IN_0_42(20) => 
        \DATA_OUT_0_42[20]\, DATA_IN_0_42(19) => 
        \DATA_OUT_0_42[19]\, DATA_IN_0_42(18) => 
        \DATA_OUT_0_42[18]\, DATA_IN_0_42(17) => 
        \DATA_OUT_0_42[17]\, DATA_IN_0_42(16) => 
        \DATA_OUT_0_42[16]\, DATA_IN_0_42(15) => 
        \DATA_OUT_0_42[15]\, DATA_IN_0_42(14) => 
        \DATA_OUT_0_42[14]\, DATA_IN_0_42(13) => 
        \DATA_OUT_0_42[13]\, DATA_IN_0_42(12) => 
        \DATA_OUT_0_42[12]\, DATA_IN_0_42(11) => 
        \DATA_OUT_0_42[11]\, DATA_IN_0_42(10) => 
        \DATA_OUT_0_42[10]\, DATA_IN_0_42(9) => 
        \DATA_OUT_0_42[9]\, DATA_IN_0_42(8) => \DATA_OUT_0_42[8]\, 
        DATA_IN_0_42(7) => \DATA_OUT_0_42[7]\, DATA_IN_0_42(6)
         => \DATA_OUT_0_42[6]\, DATA_IN_0_42(5) => 
        \DATA_OUT_0_42[5]\, DATA_IN_0_42(4) => \DATA_OUT_0_42[4]\, 
        DATA_IN_0_42(3) => \DATA_OUT_0_42[3]\, DATA_IN_0_42(2)
         => \DATA_OUT_0_42[2]\, DATA_IN_0_42(1) => 
        \DATA_OUT_0_42[1]\, DATA_IN_0_42(0) => \DATA_OUT_0_42[0]\, 
        DATA_IN_0_43(25) => \DATA_OUT_0_43[25]\, DATA_IN_0_43(24)
         => \DATA_OUT_0_43[24]\, DATA_IN_0_43(23) => 
        \DATA_OUT_0_43[23]\, DATA_IN_0_43(22) => 
        \DATA_OUT_0_43[22]\, DATA_IN_0_43(21) => 
        \DATA_OUT_0_43[21]\, DATA_IN_0_43(20) => 
        \DATA_OUT_0_43[20]\, DATA_IN_0_43(19) => 
        \DATA_OUT_0_43[19]\, DATA_IN_0_43(18) => 
        \DATA_OUT_0_43[18]\, DATA_IN_0_43(17) => 
        \DATA_OUT_0_43[17]\, DATA_IN_0_43(16) => 
        \DATA_OUT_0_43[16]\, DATA_IN_0_43(15) => 
        \DATA_OUT_0_43[15]\, DATA_IN_0_43(14) => 
        \DATA_OUT_0_43[14]\, DATA_IN_0_43(13) => 
        \DATA_OUT_0_43[13]\, DATA_IN_0_43(12) => 
        \DATA_OUT_0_43[12]\, DATA_IN_0_43(11) => 
        \DATA_OUT_0_43[11]\, DATA_IN_0_43(10) => 
        \DATA_OUT_0_43[10]\, DATA_IN_0_43(9) => 
        \DATA_OUT_0_43[9]\, DATA_IN_0_43(8) => \DATA_OUT_0_43[8]\, 
        DATA_IN_0_43(7) => \DATA_OUT_0_43[7]\, DATA_IN_0_43(6)
         => \DATA_OUT_0_43[6]\, DATA_IN_0_43(5) => 
        \DATA_OUT_0_43[5]\, DATA_IN_0_43(4) => \DATA_OUT_0_43[4]\, 
        DATA_IN_0_43(3) => \DATA_OUT_0_43[3]\, DATA_IN_0_43(2)
         => \DATA_OUT_0_43[2]\, DATA_IN_0_43(1) => 
        \DATA_OUT_0_43[1]\, DATA_IN_0_43(0) => \DATA_OUT_0_43[0]\, 
        DATA_IN_0_44(25) => \DATA_OUT_0_44[25]\, DATA_IN_0_44(24)
         => \DATA_OUT_0_44[24]\, DATA_IN_0_44(23) => 
        \DATA_OUT_0_44[23]\, DATA_IN_0_44(22) => 
        \DATA_OUT_0_44[22]\, DATA_IN_0_44(21) => 
        \DATA_OUT_0_44[21]\, DATA_IN_0_44(20) => 
        \DATA_OUT_0_44[20]\, DATA_IN_0_44(19) => 
        \DATA_OUT_0_44[19]\, DATA_IN_0_44(18) => 
        \DATA_OUT_0_44[18]\, DATA_IN_0_44(17) => 
        \DATA_OUT_0_44[17]\, DATA_IN_0_44(16) => 
        \DATA_OUT_0_44[16]\, DATA_IN_0_44(15) => 
        \DATA_OUT_0_44[15]\, DATA_IN_0_44(14) => 
        \DATA_OUT_0_44[14]\, DATA_IN_0_44(13) => 
        \DATA_OUT_0_44[13]\, DATA_IN_0_44(12) => 
        \DATA_OUT_0_44[12]\, DATA_IN_0_44(11) => 
        \DATA_OUT_0_44[11]\, DATA_IN_0_44(10) => 
        \DATA_OUT_0_44[10]\, DATA_IN_0_44(9) => 
        \DATA_OUT_0_44[9]\, DATA_IN_0_44(8) => \DATA_OUT_0_44[8]\, 
        DATA_IN_0_44(7) => \DATA_OUT_0_44[7]\, DATA_IN_0_44(6)
         => \DATA_OUT_0_44[6]\, DATA_IN_0_44(5) => 
        \DATA_OUT_0_44[5]\, DATA_IN_0_44(4) => \DATA_OUT_0_44[4]\, 
        DATA_IN_0_44(3) => \DATA_OUT_0_44[3]\, DATA_IN_0_44(2)
         => \DATA_OUT_0_44[2]\, DATA_IN_0_44(1) => 
        \DATA_OUT_0_44[1]\, DATA_IN_0_44(0) => \DATA_OUT_0_44[0]\, 
        DATA_IN_0_45(25) => \DATA_OUT_0_45[25]\, DATA_IN_0_45(24)
         => \DATA_OUT_0_45[24]\, DATA_IN_0_45(23) => 
        \DATA_OUT_0_45[23]\, DATA_IN_0_45(22) => 
        \DATA_OUT_0_45[22]\, DATA_IN_0_45(21) => 
        \DATA_OUT_0_45[21]\, DATA_IN_0_45(20) => 
        \DATA_OUT_0_45[20]\, DATA_IN_0_45(19) => 
        \DATA_OUT_0_45[19]\, DATA_IN_0_45(18) => 
        \DATA_OUT_0_45[18]\, DATA_IN_0_45(17) => 
        \DATA_OUT_0_45[17]\, DATA_IN_0_45(16) => 
        \DATA_OUT_0_45[16]\, DATA_IN_0_45(15) => 
        \DATA_OUT_0_45[15]\, DATA_IN_0_45(14) => 
        \DATA_OUT_0_45[14]\, DATA_IN_0_45(13) => 
        \DATA_OUT_0_45[13]\, DATA_IN_0_45(12) => 
        \DATA_OUT_0_45[12]\, DATA_IN_0_45(11) => 
        \DATA_OUT_0_45[11]\, DATA_IN_0_45(10) => 
        \DATA_OUT_0_45[10]\, DATA_IN_0_45(9) => 
        \DATA_OUT_0_45[9]\, DATA_IN_0_45(8) => \DATA_OUT_0_45[8]\, 
        DATA_IN_0_45(7) => \DATA_OUT_0_45[7]\, DATA_IN_0_45(6)
         => \DATA_OUT_0_45[6]\, DATA_IN_0_45(5) => 
        \DATA_OUT_0_45[5]\, DATA_IN_0_45(4) => \DATA_OUT_0_45[4]\, 
        DATA_IN_0_45(3) => \DATA_OUT_0_45[3]\, DATA_IN_0_45(2)
         => \DATA_OUT_0_45[2]\, DATA_IN_0_45(1) => 
        \DATA_OUT_0_45[1]\, DATA_IN_0_45(0) => \DATA_OUT_0_45[0]\, 
        DATA_IN_0_46(25) => \DATA_OUT_0_46[25]\, DATA_IN_0_46(24)
         => \DATA_OUT_0_46[24]\, DATA_IN_0_46(23) => 
        \DATA_OUT_0_46[23]\, DATA_IN_0_46(22) => 
        \DATA_OUT_0_46[22]\, DATA_IN_0_46(21) => 
        \DATA_OUT_0_46[21]\, DATA_IN_0_46(20) => 
        \DATA_OUT_0_46[20]\, DATA_IN_0_46(19) => 
        \DATA_OUT_0_46[19]\, DATA_IN_0_46(18) => 
        \DATA_OUT_0_46[18]\, DATA_IN_0_46(17) => 
        \DATA_OUT_0_46[17]\, DATA_IN_0_46(16) => 
        \DATA_OUT_0_46[16]\, DATA_IN_0_46(15) => 
        \DATA_OUT_0_46[15]\, DATA_IN_0_46(14) => 
        \DATA_OUT_0_46[14]\, DATA_IN_0_46(13) => 
        \DATA_OUT_0_46[13]\, DATA_IN_0_46(12) => 
        \DATA_OUT_0_46[12]\, DATA_IN_0_46(11) => 
        \DATA_OUT_0_46[11]\, DATA_IN_0_46(10) => 
        \DATA_OUT_0_46[10]\, DATA_IN_0_46(9) => 
        \DATA_OUT_0_46[9]\, DATA_IN_0_46(8) => \DATA_OUT_0_46[8]\, 
        DATA_IN_0_46(7) => \DATA_OUT_0_46[7]\, DATA_IN_0_46(6)
         => \DATA_OUT_0_46[6]\, DATA_IN_0_46(5) => 
        \DATA_OUT_0_46[5]\, DATA_IN_0_46(4) => \DATA_OUT_0_46[4]\, 
        DATA_IN_0_46(3) => \DATA_OUT_0_46[3]\, DATA_IN_0_46(2)
         => \DATA_OUT_0_46[2]\, DATA_IN_0_46(1) => 
        \DATA_OUT_0_46[1]\, DATA_IN_0_46(0) => \DATA_OUT_0_46[0]\, 
        DATA_IN_0_47(25) => \DATA_OUT_0_47[25]\, DATA_IN_0_47(24)
         => \DATA_OUT_0_47[24]\, DATA_IN_0_47(23) => 
        \DATA_OUT_0_47[23]\, DATA_IN_0_47(22) => 
        \DATA_OUT_0_47[22]\, DATA_IN_0_47(21) => 
        \DATA_OUT_0_47[21]\, DATA_IN_0_47(20) => 
        \DATA_OUT_0_47[20]\, DATA_IN_0_47(19) => 
        \DATA_OUT_0_47[19]\, DATA_IN_0_47(18) => 
        \DATA_OUT_0_47[18]\, DATA_IN_0_47(17) => 
        \DATA_OUT_0_47[17]\, DATA_IN_0_47(16) => 
        \DATA_OUT_0_47[16]\, DATA_IN_0_47(15) => 
        \DATA_OUT_0_47[15]\, DATA_IN_0_47(14) => 
        \DATA_OUT_0_47[14]\, DATA_IN_0_47(13) => 
        \DATA_OUT_0_47[13]\, DATA_IN_0_47(12) => 
        \DATA_OUT_0_47[12]\, DATA_IN_0_47(11) => 
        \DATA_OUT_0_47[11]\, DATA_IN_0_47(10) => 
        \DATA_OUT_0_47[10]\, DATA_IN_0_47(9) => 
        \DATA_OUT_0_47[9]\, DATA_IN_0_47(8) => \DATA_OUT_0_47[8]\, 
        DATA_IN_0_47(7) => \DATA_OUT_0_47[7]\, DATA_IN_0_47(6)
         => \DATA_OUT_0_47[6]\, DATA_IN_0_47(5) => 
        \DATA_OUT_0_47[5]\, DATA_IN_0_47(4) => \DATA_OUT_0_47[4]\, 
        DATA_IN_0_47(3) => \DATA_OUT_0_47[3]\, DATA_IN_0_47(2)
         => \DATA_OUT_0_47[2]\, DATA_IN_0_47(1) => 
        \DATA_OUT_0_47[1]\, DATA_IN_0_47(0) => \DATA_OUT_0_47[0]\, 
        DATA_IN_0_48(25) => \DATA_OUT_0_48[25]\, DATA_IN_0_48(24)
         => \DATA_OUT_0_48[24]\, DATA_IN_0_48(23) => 
        \DATA_OUT_0_48[23]\, DATA_IN_0_48(22) => 
        \DATA_OUT_0_48[22]\, DATA_IN_0_48(21) => 
        \DATA_OUT_0_48[21]\, DATA_IN_0_48(20) => 
        \DATA_OUT_0_48[20]\, DATA_IN_0_48(19) => 
        \DATA_OUT_0_48[19]\, DATA_IN_0_48(18) => 
        \DATA_OUT_0_48[18]\, DATA_IN_0_48(17) => 
        \DATA_OUT_0_48[17]\, DATA_IN_0_48(16) => 
        \DATA_OUT_0_48[16]\, DATA_IN_0_48(15) => 
        \DATA_OUT_0_48[15]\, DATA_IN_0_48(14) => 
        \DATA_OUT_0_48[14]\, DATA_IN_0_48(13) => 
        \DATA_OUT_0_48[13]\, DATA_IN_0_48(12) => 
        \DATA_OUT_0_48[12]\, DATA_IN_0_48(11) => 
        \DATA_OUT_0_48[11]\, DATA_IN_0_48(10) => 
        \DATA_OUT_0_48[10]\, DATA_IN_0_48(9) => 
        \DATA_OUT_0_48[9]\, DATA_IN_0_48(8) => \DATA_OUT_0_48[8]\, 
        DATA_IN_0_48(7) => \DATA_OUT_0_48[7]\, DATA_IN_0_48(6)
         => \DATA_OUT_0_48[6]\, DATA_IN_0_48(5) => 
        \DATA_OUT_0_48[5]\, DATA_IN_0_48(4) => \DATA_OUT_0_48[4]\, 
        DATA_IN_0_48(3) => \DATA_OUT_0_48[3]\, DATA_IN_0_48(2)
         => \DATA_OUT_0_48[2]\, DATA_IN_0_48(1) => 
        \DATA_OUT_0_48[1]\, DATA_IN_0_48(0) => \DATA_OUT_0_48[0]\, 
        DATA_IN_0_49(25) => \DATA_OUT_0_49[25]\, DATA_IN_0_49(24)
         => \DATA_OUT_0_49[24]\, DATA_IN_0_49(23) => 
        \DATA_OUT_0_49[23]\, DATA_IN_0_49(22) => 
        \DATA_OUT_0_49[22]\, DATA_IN_0_49(21) => 
        \DATA_OUT_0_49[21]\, DATA_IN_0_49(20) => 
        \DATA_OUT_0_49[20]\, DATA_IN_0_49(19) => 
        \DATA_OUT_0_49[19]\, DATA_IN_0_49(18) => 
        \DATA_OUT_0_49[18]\, DATA_IN_0_49(17) => 
        \DATA_OUT_0_49[17]\, DATA_IN_0_49(16) => 
        \DATA_OUT_0_49[16]\, DATA_IN_0_49(15) => 
        \DATA_OUT_0_49[15]\, DATA_IN_0_49(14) => 
        \DATA_OUT_0_49[14]\, DATA_IN_0_49(13) => 
        \DATA_OUT_0_49[13]\, DATA_IN_0_49(12) => 
        \DATA_OUT_0_49[12]\, DATA_IN_0_49(11) => 
        \DATA_OUT_0_49[11]\, DATA_IN_0_49(10) => 
        \DATA_OUT_0_49[10]\, DATA_IN_0_49(9) => 
        \DATA_OUT_0_49[9]\, DATA_IN_0_49(8) => \DATA_OUT_0_49[8]\, 
        DATA_IN_0_49(7) => \DATA_OUT_0_49[7]\, DATA_IN_0_49(6)
         => \DATA_OUT_0_49[6]\, DATA_IN_0_49(5) => 
        \DATA_OUT_0_49[5]\, DATA_IN_0_49(4) => \DATA_OUT_0_49[4]\, 
        DATA_IN_0_49(3) => \DATA_OUT_0_49[3]\, DATA_IN_0_49(2)
         => \DATA_OUT_0_49[2]\, DATA_IN_0_49(1) => 
        \DATA_OUT_0_49[1]\, DATA_IN_0_49(0) => \DATA_OUT_0_49[0]\, 
        DATA_IN_0_50(25) => \DATA_OUT_0_50[25]\, DATA_IN_0_50(24)
         => \DATA_OUT_0_50[24]\, DATA_IN_0_50(23) => 
        \DATA_OUT_0_50[23]\, DATA_IN_0_50(22) => 
        \DATA_OUT_0_50[22]\, DATA_IN_0_50(21) => 
        \DATA_OUT_0_50[21]\, DATA_IN_0_50(20) => 
        \DATA_OUT_0_50[20]\, DATA_IN_0_50(19) => 
        \DATA_OUT_0_50[19]\, DATA_IN_0_50(18) => 
        \DATA_OUT_0_50[18]\, DATA_IN_0_50(17) => 
        \DATA_OUT_0_50[17]\, DATA_IN_0_50(16) => 
        \DATA_OUT_0_50[16]\, DATA_IN_0_50(15) => 
        \DATA_OUT_0_50[15]\, DATA_IN_0_50(14) => 
        \DATA_OUT_0_50[14]\, DATA_IN_0_50(13) => 
        \DATA_OUT_0_50[13]\, DATA_IN_0_50(12) => 
        \DATA_OUT_0_50[12]\, DATA_IN_0_50(11) => 
        \DATA_OUT_0_50[11]\, DATA_IN_0_50(10) => 
        \DATA_OUT_0_50[10]\, DATA_IN_0_50(9) => 
        \DATA_OUT_0_50[9]\, DATA_IN_0_50(8) => \DATA_OUT_0_50[8]\, 
        DATA_IN_0_50(7) => \DATA_OUT_0_50[7]\, DATA_IN_0_50(6)
         => \DATA_OUT_0_50[6]\, DATA_IN_0_50(5) => 
        \DATA_OUT_0_50[5]\, DATA_IN_0_50(4) => \DATA_OUT_0_50[4]\, 
        DATA_IN_0_50(3) => \DATA_OUT_0_50[3]\, DATA_IN_0_50(2)
         => \DATA_OUT_0_50[2]\, DATA_IN_0_50(1) => 
        \DATA_OUT_0_50[1]\, DATA_IN_0_50(0) => \DATA_OUT_0_50[0]\, 
        DATA_IN_0_51(25) => \DATA_OUT_0_51[25]\, DATA_IN_0_51(24)
         => \DATA_OUT_0_51[24]\, DATA_IN_0_51(23) => 
        \DATA_OUT_0_51[23]\, DATA_IN_0_51(22) => 
        \DATA_OUT_0_51[22]\, DATA_IN_0_51(21) => 
        \DATA_OUT_0_51[21]\, DATA_IN_0_51(20) => 
        \DATA_OUT_0_51[20]\, DATA_IN_0_51(19) => 
        \DATA_OUT_0_51[19]\, DATA_IN_0_51(18) => 
        \DATA_OUT_0_51[18]\, DATA_IN_0_51(17) => 
        \DATA_OUT_0_51[17]\, DATA_IN_0_51(16) => 
        \DATA_OUT_0_51[16]\, DATA_IN_0_51(15) => 
        \DATA_OUT_0_51[15]\, DATA_IN_0_51(14) => 
        \DATA_OUT_0_51[14]\, DATA_IN_0_51(13) => 
        \DATA_OUT_0_51[13]\, DATA_IN_0_51(12) => 
        \DATA_OUT_0_51[12]\, DATA_IN_0_51(11) => 
        \DATA_OUT_0_51[11]\, DATA_IN_0_51(10) => 
        \DATA_OUT_0_51[10]\, DATA_IN_0_51(9) => 
        \DATA_OUT_0_51[9]\, DATA_IN_0_51(8) => \DATA_OUT_0_51[8]\, 
        DATA_IN_0_51(7) => \DATA_OUT_0_51[7]\, DATA_IN_0_51(6)
         => \DATA_OUT_0_51[6]\, DATA_IN_0_51(5) => 
        \DATA_OUT_0_51[5]\, DATA_IN_0_51(4) => \DATA_OUT_0_51[4]\, 
        DATA_IN_0_51(3) => \DATA_OUT_0_51[3]\, DATA_IN_0_51(2)
         => \DATA_OUT_0_51[2]\, DATA_IN_0_51(1) => 
        \DATA_OUT_0_51[1]\, DATA_IN_0_51(0) => \DATA_OUT_0_51[0]\, 
        DATA_IN_1_0(25) => \DATA_OUT_1_0[25]\, DATA_IN_1_0(24)
         => \DATA_OUT_1_0[24]\, DATA_IN_1_0(23) => 
        \DATA_OUT_1_0[23]\, DATA_IN_1_0(22) => \DATA_OUT_1_0[22]\, 
        DATA_IN_1_0(21) => \DATA_OUT_1_0[21]\, DATA_IN_1_0(20)
         => \DATA_OUT_1_0[20]\, DATA_IN_1_0(19) => 
        \DATA_OUT_1_0[19]\, DATA_IN_1_0(18) => \DATA_OUT_1_0[18]\, 
        DATA_IN_1_0(17) => \DATA_OUT_1_0[17]\, DATA_IN_1_0(16)
         => \DATA_OUT_1_0[16]\, DATA_IN_1_0(15) => 
        \DATA_OUT_1_0[15]\, DATA_IN_1_0(14) => \DATA_OUT_1_0[14]\, 
        DATA_IN_1_0(13) => \DATA_OUT_1_0[13]\, DATA_IN_1_0(12)
         => \DATA_OUT_1_0[12]\, DATA_IN_1_0(11) => 
        \DATA_OUT_1_0[11]\, DATA_IN_1_0(10) => \DATA_OUT_1_0[10]\, 
        DATA_IN_1_0(9) => \DATA_OUT_1_0[9]\, DATA_IN_1_0(8) => 
        \DATA_OUT_1_0[8]\, DATA_IN_1_0(7) => \DATA_OUT_1_0[7]\, 
        DATA_IN_1_0(6) => \DATA_OUT_1_0[6]\, DATA_IN_1_0(5) => 
        \DATA_OUT_1_0[5]\, DATA_IN_1_0(4) => \DATA_OUT_1_0[4]\, 
        DATA_IN_1_0(3) => \DATA_OUT_1_0[3]\, DATA_IN_1_0(2) => 
        \DATA_OUT_1_0[2]\, DATA_IN_1_0(1) => \DATA_OUT_1_0[1]\, 
        DATA_IN_1_0(0) => \DATA_OUT_1_0[0]\, DATA_IN_1_1(25) => 
        \DATA_OUT_1_1[25]\, DATA_IN_1_1(24) => \DATA_OUT_1_1[24]\, 
        DATA_IN_1_1(23) => \DATA_OUT_1_1[23]\, DATA_IN_1_1(22)
         => \DATA_OUT_1_1[22]\, DATA_IN_1_1(21) => 
        \DATA_OUT_1_1[21]\, DATA_IN_1_1(20) => \DATA_OUT_1_1[20]\, 
        DATA_IN_1_1(19) => \DATA_OUT_1_1[19]\, DATA_IN_1_1(18)
         => \DATA_OUT_1_1[18]\, DATA_IN_1_1(17) => 
        \DATA_OUT_1_1[17]\, DATA_IN_1_1(16) => \DATA_OUT_1_1[16]\, 
        DATA_IN_1_1(15) => \DATA_OUT_1_1[15]\, DATA_IN_1_1(14)
         => \DATA_OUT_1_1[14]\, DATA_IN_1_1(13) => 
        \DATA_OUT_1_1[13]\, DATA_IN_1_1(12) => \DATA_OUT_1_1[12]\, 
        DATA_IN_1_1(11) => \DATA_OUT_1_1[11]\, DATA_IN_1_1(10)
         => \DATA_OUT_1_1[10]\, DATA_IN_1_1(9) => 
        \DATA_OUT_1_1[9]\, DATA_IN_1_1(8) => \DATA_OUT_1_1[8]\, 
        DATA_IN_1_1(7) => \DATA_OUT_1_1[7]\, DATA_IN_1_1(6) => 
        \DATA_OUT_1_1[6]\, DATA_IN_1_1(5) => \DATA_OUT_1_1[5]\, 
        DATA_IN_1_1(4) => \DATA_OUT_1_1[4]\, DATA_IN_1_1(3) => 
        \DATA_OUT_1_1[3]\, DATA_IN_1_1(2) => \DATA_OUT_1_1[2]\, 
        DATA_IN_1_1(1) => \DATA_OUT_1_1[1]\, DATA_IN_1_1(0) => 
        \DATA_OUT_1_1[0]\, DATA_IN_1_2(25) => \DATA_OUT_1_2[25]\, 
        DATA_IN_1_2(24) => \DATA_OUT_1_2[24]\, DATA_IN_1_2(23)
         => \DATA_OUT_1_2[23]\, DATA_IN_1_2(22) => 
        \DATA_OUT_1_2[22]\, DATA_IN_1_2(21) => \DATA_OUT_1_2[21]\, 
        DATA_IN_1_2(20) => \DATA_OUT_1_2[20]\, DATA_IN_1_2(19)
         => \DATA_OUT_1_2[19]\, DATA_IN_1_2(18) => 
        \DATA_OUT_1_2[18]\, DATA_IN_1_2(17) => \DATA_OUT_1_2[17]\, 
        DATA_IN_1_2(16) => \DATA_OUT_1_2[16]\, DATA_IN_1_2(15)
         => \DATA_OUT_1_2[15]\, DATA_IN_1_2(14) => 
        \DATA_OUT_1_2[14]\, DATA_IN_1_2(13) => \DATA_OUT_1_2[13]\, 
        DATA_IN_1_2(12) => \DATA_OUT_1_2[12]\, DATA_IN_1_2(11)
         => \DATA_OUT_1_2[11]\, DATA_IN_1_2(10) => 
        \DATA_OUT_1_2[10]\, DATA_IN_1_2(9) => \DATA_OUT_1_2[9]\, 
        DATA_IN_1_2(8) => \DATA_OUT_1_2[8]\, DATA_IN_1_2(7) => 
        \DATA_OUT_1_2[7]\, DATA_IN_1_2(6) => \DATA_OUT_1_2[6]\, 
        DATA_IN_1_2(5) => \DATA_OUT_1_2[5]\, DATA_IN_1_2(4) => 
        \DATA_OUT_1_2[4]\, DATA_IN_1_2(3) => \DATA_OUT_1_2[3]\, 
        DATA_IN_1_2(2) => \DATA_OUT_1_2[2]\, DATA_IN_1_2(1) => 
        \DATA_OUT_1_2[1]\, DATA_IN_1_2(0) => \DATA_OUT_1_2[0]\, 
        DATA_IN_1_3(25) => \DATA_OUT_1_3[25]\, DATA_IN_1_3(24)
         => \DATA_OUT_1_3[24]\, DATA_IN_1_3(23) => 
        \DATA_OUT_1_3[23]\, DATA_IN_1_3(22) => \DATA_OUT_1_3[22]\, 
        DATA_IN_1_3(21) => \DATA_OUT_1_3[21]\, DATA_IN_1_3(20)
         => \DATA_OUT_1_3[20]\, DATA_IN_1_3(19) => 
        \DATA_OUT_1_3[19]\, DATA_IN_1_3(18) => \DATA_OUT_1_3[18]\, 
        DATA_IN_1_3(17) => \DATA_OUT_1_3[17]\, DATA_IN_1_3(16)
         => \DATA_OUT_1_3[16]\, DATA_IN_1_3(15) => 
        \DATA_OUT_1_3[15]\, DATA_IN_1_3(14) => \DATA_OUT_1_3[14]\, 
        DATA_IN_1_3(13) => \DATA_OUT_1_3[13]\, DATA_IN_1_3(12)
         => \DATA_OUT_1_3[12]\, DATA_IN_1_3(11) => 
        \DATA_OUT_1_3[11]\, DATA_IN_1_3(10) => \DATA_OUT_1_3[10]\, 
        DATA_IN_1_3(9) => \DATA_OUT_1_3[9]\, DATA_IN_1_3(8) => 
        \DATA_OUT_1_3[8]\, DATA_IN_1_3(7) => \DATA_OUT_1_3[7]\, 
        DATA_IN_1_3(6) => \DATA_OUT_1_3[6]\, DATA_IN_1_3(5) => 
        \DATA_OUT_1_3[5]\, DATA_IN_1_3(4) => \DATA_OUT_1_3[4]\, 
        DATA_IN_1_3(3) => \DATA_OUT_1_3[3]\, DATA_IN_1_3(2) => 
        \DATA_OUT_1_3[2]\, DATA_IN_1_3(1) => \DATA_OUT_1_3[1]\, 
        DATA_IN_1_3(0) => \DATA_OUT_1_3[0]\, DATA_IN_1_4(25) => 
        \DATA_OUT_1_4[25]\, DATA_IN_1_4(24) => \DATA_OUT_1_4[24]\, 
        DATA_IN_1_4(23) => \DATA_OUT_1_4[23]\, DATA_IN_1_4(22)
         => \DATA_OUT_1_4[22]\, DATA_IN_1_4(21) => 
        \DATA_OUT_1_4[21]\, DATA_IN_1_4(20) => \DATA_OUT_1_4[20]\, 
        DATA_IN_1_4(19) => \DATA_OUT_1_4[19]\, DATA_IN_1_4(18)
         => \DATA_OUT_1_4[18]\, DATA_IN_1_4(17) => 
        \DATA_OUT_1_4[17]\, DATA_IN_1_4(16) => \DATA_OUT_1_4[16]\, 
        DATA_IN_1_4(15) => \DATA_OUT_1_4[15]\, DATA_IN_1_4(14)
         => \DATA_OUT_1_4[14]\, DATA_IN_1_4(13) => 
        \DATA_OUT_1_4[13]\, DATA_IN_1_4(12) => \DATA_OUT_1_4[12]\, 
        DATA_IN_1_4(11) => \DATA_OUT_1_4[11]\, DATA_IN_1_4(10)
         => \DATA_OUT_1_4[10]\, DATA_IN_1_4(9) => 
        \DATA_OUT_1_4[9]\, DATA_IN_1_4(8) => \DATA_OUT_1_4[8]\, 
        DATA_IN_1_4(7) => \DATA_OUT_1_4[7]\, DATA_IN_1_4(6) => 
        \DATA_OUT_1_4[6]\, DATA_IN_1_4(5) => \DATA_OUT_1_4[5]\, 
        DATA_IN_1_4(4) => \DATA_OUT_1_4[4]\, DATA_IN_1_4(3) => 
        \DATA_OUT_1_4[3]\, DATA_IN_1_4(2) => \DATA_OUT_1_4[2]\, 
        DATA_IN_1_4(1) => \DATA_OUT_1_4[1]\, DATA_IN_1_4(0) => 
        \DATA_OUT_1_4[0]\, DATA_IN_1_5(25) => \DATA_OUT_1_5[25]\, 
        DATA_IN_1_5(24) => \DATA_OUT_1_5[24]\, DATA_IN_1_5(23)
         => \DATA_OUT_1_5[23]\, DATA_IN_1_5(22) => 
        \DATA_OUT_1_5[22]\, DATA_IN_1_5(21) => \DATA_OUT_1_5[21]\, 
        DATA_IN_1_5(20) => \DATA_OUT_1_5[20]\, DATA_IN_1_5(19)
         => \DATA_OUT_1_5[19]\, DATA_IN_1_5(18) => 
        \DATA_OUT_1_5[18]\, DATA_IN_1_5(17) => \DATA_OUT_1_5[17]\, 
        DATA_IN_1_5(16) => \DATA_OUT_1_5[16]\, DATA_IN_1_5(15)
         => \DATA_OUT_1_5[15]\, DATA_IN_1_5(14) => 
        \DATA_OUT_1_5[14]\, DATA_IN_1_5(13) => \DATA_OUT_1_5[13]\, 
        DATA_IN_1_5(12) => \DATA_OUT_1_5[12]\, DATA_IN_1_5(11)
         => \DATA_OUT_1_5[11]\, DATA_IN_1_5(10) => 
        \DATA_OUT_1_5[10]\, DATA_IN_1_5(9) => \DATA_OUT_1_5[9]\, 
        DATA_IN_1_5(8) => \DATA_OUT_1_5[8]\, DATA_IN_1_5(7) => 
        \DATA_OUT_1_5[7]\, DATA_IN_1_5(6) => \DATA_OUT_1_5[6]\, 
        DATA_IN_1_5(5) => \DATA_OUT_1_5[5]\, DATA_IN_1_5(4) => 
        \DATA_OUT_1_5[4]\, DATA_IN_1_5(3) => \DATA_OUT_1_5[3]\, 
        DATA_IN_1_5(2) => \DATA_OUT_1_5[2]\, DATA_IN_1_5(1) => 
        \DATA_OUT_1_5[1]\, DATA_IN_1_5(0) => \DATA_OUT_1_5[0]\, 
        DATA_IN_1_6(25) => \DATA_OUT_1_6[25]\, DATA_IN_1_6(24)
         => \DATA_OUT_1_6[24]\, DATA_IN_1_6(23) => 
        \DATA_OUT_1_6[23]\, DATA_IN_1_6(22) => \DATA_OUT_1_6[22]\, 
        DATA_IN_1_6(21) => \DATA_OUT_1_6[21]\, DATA_IN_1_6(20)
         => \DATA_OUT_1_6[20]\, DATA_IN_1_6(19) => 
        \DATA_OUT_1_6[19]\, DATA_IN_1_6(18) => \DATA_OUT_1_6[18]\, 
        DATA_IN_1_6(17) => \DATA_OUT_1_6[17]\, DATA_IN_1_6(16)
         => \DATA_OUT_1_6[16]\, DATA_IN_1_6(15) => 
        \DATA_OUT_1_6[15]\, DATA_IN_1_6(14) => \DATA_OUT_1_6[14]\, 
        DATA_IN_1_6(13) => \DATA_OUT_1_6[13]\, DATA_IN_1_6(12)
         => \DATA_OUT_1_6[12]\, DATA_IN_1_6(11) => 
        \DATA_OUT_1_6[11]\, DATA_IN_1_6(10) => \DATA_OUT_1_6[10]\, 
        DATA_IN_1_6(9) => \DATA_OUT_1_6[9]\, DATA_IN_1_6(8) => 
        \DATA_OUT_1_6[8]\, DATA_IN_1_6(7) => \DATA_OUT_1_6[7]\, 
        DATA_IN_1_6(6) => \DATA_OUT_1_6[6]\, DATA_IN_1_6(5) => 
        \DATA_OUT_1_6[5]\, DATA_IN_1_6(4) => \DATA_OUT_1_6[4]\, 
        DATA_IN_1_6(3) => \DATA_OUT_1_6[3]\, DATA_IN_1_6(2) => 
        \DATA_OUT_1_6[2]\, DATA_IN_1_6(1) => \DATA_OUT_1_6[1]\, 
        DATA_IN_1_6(0) => \DATA_OUT_1_6[0]\, DATA_IN_1_7(25) => 
        \DATA_OUT_1_7[25]\, DATA_IN_1_7(24) => \DATA_OUT_1_7[24]\, 
        DATA_IN_1_7(23) => \DATA_OUT_1_7[23]\, DATA_IN_1_7(22)
         => \DATA_OUT_1_7[22]\, DATA_IN_1_7(21) => 
        \DATA_OUT_1_7[21]\, DATA_IN_1_7(20) => \DATA_OUT_1_7[20]\, 
        DATA_IN_1_7(19) => \DATA_OUT_1_7[19]\, DATA_IN_1_7(18)
         => \DATA_OUT_1_7[18]\, DATA_IN_1_7(17) => 
        \DATA_OUT_1_7[17]\, DATA_IN_1_7(16) => \DATA_OUT_1_7[16]\, 
        DATA_IN_1_7(15) => \DATA_OUT_1_7[15]\, DATA_IN_1_7(14)
         => \DATA_OUT_1_7[14]\, DATA_IN_1_7(13) => 
        \DATA_OUT_1_7[13]\, DATA_IN_1_7(12) => \DATA_OUT_1_7[12]\, 
        DATA_IN_1_7(11) => \DATA_OUT_1_7[11]\, DATA_IN_1_7(10)
         => \DATA_OUT_1_7[10]\, DATA_IN_1_7(9) => 
        \DATA_OUT_1_7[9]\, DATA_IN_1_7(8) => \DATA_OUT_1_7[8]\, 
        DATA_IN_1_7(7) => \DATA_OUT_1_7[7]\, DATA_IN_1_7(6) => 
        \DATA_OUT_1_7[6]\, DATA_IN_1_7(5) => \DATA_OUT_1_7[5]\, 
        DATA_IN_1_7(4) => \DATA_OUT_1_7[4]\, DATA_IN_1_7(3) => 
        \DATA_OUT_1_7[3]\, DATA_IN_1_7(2) => \DATA_OUT_1_7[2]\, 
        DATA_IN_1_7(1) => \DATA_OUT_1_7[1]\, DATA_IN_1_7(0) => 
        \DATA_OUT_1_7[0]\, DATA_IN_1_8(25) => \DATA_OUT_1_8[25]\, 
        DATA_IN_1_8(24) => \DATA_OUT_1_8[24]\, DATA_IN_1_8(23)
         => \DATA_OUT_1_8[23]\, DATA_IN_1_8(22) => 
        \DATA_OUT_1_8[22]\, DATA_IN_1_8(21) => \DATA_OUT_1_8[21]\, 
        DATA_IN_1_8(20) => \DATA_OUT_1_8[20]\, DATA_IN_1_8(19)
         => \DATA_OUT_1_8[19]\, DATA_IN_1_8(18) => 
        \DATA_OUT_1_8[18]\, DATA_IN_1_8(17) => \DATA_OUT_1_8[17]\, 
        DATA_IN_1_8(16) => \DATA_OUT_1_8[16]\, DATA_IN_1_8(15)
         => \DATA_OUT_1_8[15]\, DATA_IN_1_8(14) => 
        \DATA_OUT_1_8[14]\, DATA_IN_1_8(13) => \DATA_OUT_1_8[13]\, 
        DATA_IN_1_8(12) => \DATA_OUT_1_8[12]\, DATA_IN_1_8(11)
         => \DATA_OUT_1_8[11]\, DATA_IN_1_8(10) => 
        \DATA_OUT_1_8[10]\, DATA_IN_1_8(9) => \DATA_OUT_1_8[9]\, 
        DATA_IN_1_8(8) => \DATA_OUT_1_8[8]\, DATA_IN_1_8(7) => 
        \DATA_OUT_1_8[7]\, DATA_IN_1_8(6) => \DATA_OUT_1_8[6]\, 
        DATA_IN_1_8(5) => \DATA_OUT_1_8[5]\, DATA_IN_1_8(4) => 
        \DATA_OUT_1_8[4]\, DATA_IN_1_8(3) => \DATA_OUT_1_8[3]\, 
        DATA_IN_1_8(2) => \DATA_OUT_1_8[2]\, DATA_IN_1_8(1) => 
        \DATA_OUT_1_8[1]\, DATA_IN_1_8(0) => \DATA_OUT_1_8[0]\, 
        DATA_IN_1_9(25) => \DATA_OUT_1_9[25]\, DATA_IN_1_9(24)
         => \DATA_OUT_1_9[24]\, DATA_IN_1_9(23) => 
        \DATA_OUT_1_9[23]\, DATA_IN_1_9(22) => \DATA_OUT_1_9[22]\, 
        DATA_IN_1_9(21) => \DATA_OUT_1_9[21]\, DATA_IN_1_9(20)
         => \DATA_OUT_1_9[20]\, DATA_IN_1_9(19) => 
        \DATA_OUT_1_9[19]\, DATA_IN_1_9(18) => \DATA_OUT_1_9[18]\, 
        DATA_IN_1_9(17) => \DATA_OUT_1_9[17]\, DATA_IN_1_9(16)
         => \DATA_OUT_1_9[16]\, DATA_IN_1_9(15) => 
        \DATA_OUT_1_9[15]\, DATA_IN_1_9(14) => \DATA_OUT_1_9[14]\, 
        DATA_IN_1_9(13) => \DATA_OUT_1_9[13]\, DATA_IN_1_9(12)
         => \DATA_OUT_1_9[12]\, DATA_IN_1_9(11) => 
        \DATA_OUT_1_9[11]\, DATA_IN_1_9(10) => \DATA_OUT_1_9[10]\, 
        DATA_IN_1_9(9) => \DATA_OUT_1_9[9]\, DATA_IN_1_9(8) => 
        \DATA_OUT_1_9[8]\, DATA_IN_1_9(7) => \DATA_OUT_1_9[7]\, 
        DATA_IN_1_9(6) => \DATA_OUT_1_9[6]\, DATA_IN_1_9(5) => 
        \DATA_OUT_1_9[5]\, DATA_IN_1_9(4) => \DATA_OUT_1_9[4]\, 
        DATA_IN_1_9(3) => \DATA_OUT_1_9[3]\, DATA_IN_1_9(2) => 
        \DATA_OUT_1_9[2]\, DATA_IN_1_9(1) => \DATA_OUT_1_9[1]\, 
        DATA_IN_1_9(0) => \DATA_OUT_1_9[0]\, DATA_IN_1_10(25) => 
        \DATA_OUT_1_10[25]\, DATA_IN_1_10(24) => 
        \DATA_OUT_1_10[24]\, DATA_IN_1_10(23) => 
        \DATA_OUT_1_10[23]\, DATA_IN_1_10(22) => 
        \DATA_OUT_1_10[22]\, DATA_IN_1_10(21) => 
        \DATA_OUT_1_10[21]\, DATA_IN_1_10(20) => 
        \DATA_OUT_1_10[20]\, DATA_IN_1_10(19) => 
        \DATA_OUT_1_10[19]\, DATA_IN_1_10(18) => 
        \DATA_OUT_1_10[18]\, DATA_IN_1_10(17) => 
        \DATA_OUT_1_10[17]\, DATA_IN_1_10(16) => 
        \DATA_OUT_1_10[16]\, DATA_IN_1_10(15) => 
        \DATA_OUT_1_10[15]\, DATA_IN_1_10(14) => 
        \DATA_OUT_1_10[14]\, DATA_IN_1_10(13) => 
        \DATA_OUT_1_10[13]\, DATA_IN_1_10(12) => 
        \DATA_OUT_1_10[12]\, DATA_IN_1_10(11) => 
        \DATA_OUT_1_10[11]\, DATA_IN_1_10(10) => 
        \DATA_OUT_1_10[10]\, DATA_IN_1_10(9) => 
        \DATA_OUT_1_10[9]\, DATA_IN_1_10(8) => \DATA_OUT_1_10[8]\, 
        DATA_IN_1_10(7) => \DATA_OUT_1_10[7]\, DATA_IN_1_10(6)
         => \DATA_OUT_1_10[6]\, DATA_IN_1_10(5) => 
        \DATA_OUT_1_10[5]\, DATA_IN_1_10(4) => \DATA_OUT_1_10[4]\, 
        DATA_IN_1_10(3) => \DATA_OUT_1_10[3]\, DATA_IN_1_10(2)
         => \DATA_OUT_1_10[2]\, DATA_IN_1_10(1) => 
        \DATA_OUT_1_10[1]\, DATA_IN_1_10(0) => \DATA_OUT_1_10[0]\, 
        DATA_IN_1_11(25) => \DATA_OUT_1_11[25]\, DATA_IN_1_11(24)
         => \DATA_OUT_1_11[24]\, DATA_IN_1_11(23) => 
        \DATA_OUT_1_11[23]\, DATA_IN_1_11(22) => 
        \DATA_OUT_1_11[22]\, DATA_IN_1_11(21) => 
        \DATA_OUT_1_11[21]\, DATA_IN_1_11(20) => 
        \DATA_OUT_1_11[20]\, DATA_IN_1_11(19) => 
        \DATA_OUT_1_11[19]\, DATA_IN_1_11(18) => 
        \DATA_OUT_1_11[18]\, DATA_IN_1_11(17) => 
        \DATA_OUT_1_11[17]\, DATA_IN_1_11(16) => 
        \DATA_OUT_1_11[16]\, DATA_IN_1_11(15) => 
        \DATA_OUT_1_11[15]\, DATA_IN_1_11(14) => 
        \DATA_OUT_1_11[14]\, DATA_IN_1_11(13) => 
        \DATA_OUT_1_11[13]\, DATA_IN_1_11(12) => 
        \DATA_OUT_1_11[12]\, DATA_IN_1_11(11) => 
        \DATA_OUT_1_11[11]\, DATA_IN_1_11(10) => 
        \DATA_OUT_1_11[10]\, DATA_IN_1_11(9) => 
        \DATA_OUT_1_11[9]\, DATA_IN_1_11(8) => \DATA_OUT_1_11[8]\, 
        DATA_IN_1_11(7) => \DATA_OUT_1_11[7]\, DATA_IN_1_11(6)
         => \DATA_OUT_1_11[6]\, DATA_IN_1_11(5) => 
        \DATA_OUT_1_11[5]\, DATA_IN_1_11(4) => \DATA_OUT_1_11[4]\, 
        DATA_IN_1_11(3) => \DATA_OUT_1_11[3]\, DATA_IN_1_11(2)
         => \DATA_OUT_1_11[2]\, DATA_IN_1_11(1) => 
        \DATA_OUT_1_11[1]\, DATA_IN_1_11(0) => \DATA_OUT_1_11[0]\, 
        DATA_IN_1_12(25) => \DATA_OUT_1_12[25]\, DATA_IN_1_12(24)
         => \DATA_OUT_1_12[24]\, DATA_IN_1_12(23) => 
        \DATA_OUT_1_12[23]\, DATA_IN_1_12(22) => 
        \DATA_OUT_1_12[22]\, DATA_IN_1_12(21) => 
        \DATA_OUT_1_12[21]\, DATA_IN_1_12(20) => 
        \DATA_OUT_1_12[20]\, DATA_IN_1_12(19) => 
        \DATA_OUT_1_12[19]\, DATA_IN_1_12(18) => 
        \DATA_OUT_1_12[18]\, DATA_IN_1_12(17) => 
        \DATA_OUT_1_12[17]\, DATA_IN_1_12(16) => 
        \DATA_OUT_1_12[16]\, DATA_IN_1_12(15) => 
        \DATA_OUT_1_12[15]\, DATA_IN_1_12(14) => 
        \DATA_OUT_1_12[14]\, DATA_IN_1_12(13) => 
        \DATA_OUT_1_12[13]\, DATA_IN_1_12(12) => 
        \DATA_OUT_1_12[12]\, DATA_IN_1_12(11) => 
        \DATA_OUT_1_12[11]\, DATA_IN_1_12(10) => 
        \DATA_OUT_1_12[10]\, DATA_IN_1_12(9) => 
        \DATA_OUT_1_12[9]\, DATA_IN_1_12(8) => \DATA_OUT_1_12[8]\, 
        DATA_IN_1_12(7) => \DATA_OUT_1_12[7]\, DATA_IN_1_12(6)
         => \DATA_OUT_1_12[6]\, DATA_IN_1_12(5) => 
        \DATA_OUT_1_12[5]\, DATA_IN_1_12(4) => \DATA_OUT_1_12[4]\, 
        DATA_IN_1_12(3) => \DATA_OUT_1_12[3]\, DATA_IN_1_12(2)
         => \DATA_OUT_1_12[2]\, DATA_IN_1_12(1) => 
        \DATA_OUT_1_12[1]\, DATA_IN_1_12(0) => \DATA_OUT_1_12[0]\, 
        DATA_IN_1_13(25) => \DATA_OUT_1_13[25]\, DATA_IN_1_13(24)
         => \DATA_OUT_1_13[24]\, DATA_IN_1_13(23) => 
        \DATA_OUT_1_13[23]\, DATA_IN_1_13(22) => 
        \DATA_OUT_1_13[22]\, DATA_IN_1_13(21) => 
        \DATA_OUT_1_13[21]\, DATA_IN_1_13(20) => 
        \DATA_OUT_1_13[20]\, DATA_IN_1_13(19) => 
        \DATA_OUT_1_13[19]\, DATA_IN_1_13(18) => 
        \DATA_OUT_1_13[18]\, DATA_IN_1_13(17) => 
        \DATA_OUT_1_13[17]\, DATA_IN_1_13(16) => 
        \DATA_OUT_1_13[16]\, DATA_IN_1_13(15) => 
        \DATA_OUT_1_13[15]\, DATA_IN_1_13(14) => 
        \DATA_OUT_1_13[14]\, DATA_IN_1_13(13) => 
        \DATA_OUT_1_13[13]\, DATA_IN_1_13(12) => 
        \DATA_OUT_1_13[12]\, DATA_IN_1_13(11) => 
        \DATA_OUT_1_13[11]\, DATA_IN_1_13(10) => 
        \DATA_OUT_1_13[10]\, DATA_IN_1_13(9) => 
        \DATA_OUT_1_13[9]\, DATA_IN_1_13(8) => \DATA_OUT_1_13[8]\, 
        DATA_IN_1_13(7) => \DATA_OUT_1_13[7]\, DATA_IN_1_13(6)
         => \DATA_OUT_1_13[6]\, DATA_IN_1_13(5) => 
        \DATA_OUT_1_13[5]\, DATA_IN_1_13(4) => \DATA_OUT_1_13[4]\, 
        DATA_IN_1_13(3) => \DATA_OUT_1_13[3]\, DATA_IN_1_13(2)
         => \DATA_OUT_1_13[2]\, DATA_IN_1_13(1) => 
        \DATA_OUT_1_13[1]\, DATA_IN_1_13(0) => \DATA_OUT_1_13[0]\, 
        DATA_IN_1_14(25) => \DATA_OUT_1_14[25]\, DATA_IN_1_14(24)
         => \DATA_OUT_1_14[24]\, DATA_IN_1_14(23) => 
        \DATA_OUT_1_14[23]\, DATA_IN_1_14(22) => 
        \DATA_OUT_1_14[22]\, DATA_IN_1_14(21) => 
        \DATA_OUT_1_14[21]\, DATA_IN_1_14(20) => 
        \DATA_OUT_1_14[20]\, DATA_IN_1_14(19) => 
        \DATA_OUT_1_14[19]\, DATA_IN_1_14(18) => 
        \DATA_OUT_1_14[18]\, DATA_IN_1_14(17) => 
        \DATA_OUT_1_14[17]\, DATA_IN_1_14(16) => 
        \DATA_OUT_1_14[16]\, DATA_IN_1_14(15) => 
        \DATA_OUT_1_14[15]\, DATA_IN_1_14(14) => 
        \DATA_OUT_1_14[14]\, DATA_IN_1_14(13) => 
        \DATA_OUT_1_14[13]\, DATA_IN_1_14(12) => 
        \DATA_OUT_1_14[12]\, DATA_IN_1_14(11) => 
        \DATA_OUT_1_14[11]\, DATA_IN_1_14(10) => 
        \DATA_OUT_1_14[10]\, DATA_IN_1_14(9) => 
        \DATA_OUT_1_14[9]\, DATA_IN_1_14(8) => \DATA_OUT_1_14[8]\, 
        DATA_IN_1_14(7) => \DATA_OUT_1_14[7]\, DATA_IN_1_14(6)
         => \DATA_OUT_1_14[6]\, DATA_IN_1_14(5) => 
        \DATA_OUT_1_14[5]\, DATA_IN_1_14(4) => \DATA_OUT_1_14[4]\, 
        DATA_IN_1_14(3) => \DATA_OUT_1_14[3]\, DATA_IN_1_14(2)
         => \DATA_OUT_1_14[2]\, DATA_IN_1_14(1) => 
        \DATA_OUT_1_14[1]\, DATA_IN_1_14(0) => \DATA_OUT_1_14[0]\, 
        DATA_IN_1_15(25) => \DATA_OUT_1_15[25]\, DATA_IN_1_15(24)
         => \DATA_OUT_1_15[24]\, DATA_IN_1_15(23) => 
        \DATA_OUT_1_15[23]\, DATA_IN_1_15(22) => 
        \DATA_OUT_1_15[22]\, DATA_IN_1_15(21) => 
        \DATA_OUT_1_15[21]\, DATA_IN_1_15(20) => 
        \DATA_OUT_1_15[20]\, DATA_IN_1_15(19) => 
        \DATA_OUT_1_15[19]\, DATA_IN_1_15(18) => 
        \DATA_OUT_1_15[18]\, DATA_IN_1_15(17) => 
        \DATA_OUT_1_15[17]\, DATA_IN_1_15(16) => 
        \DATA_OUT_1_15[16]\, DATA_IN_1_15(15) => 
        \DATA_OUT_1_15[15]\, DATA_IN_1_15(14) => 
        \DATA_OUT_1_15[14]\, DATA_IN_1_15(13) => 
        \DATA_OUT_1_15[13]\, DATA_IN_1_15(12) => 
        \DATA_OUT_1_15[12]\, DATA_IN_1_15(11) => 
        \DATA_OUT_1_15[11]\, DATA_IN_1_15(10) => 
        \DATA_OUT_1_15[10]\, DATA_IN_1_15(9) => 
        \DATA_OUT_1_15[9]\, DATA_IN_1_15(8) => \DATA_OUT_1_15[8]\, 
        DATA_IN_1_15(7) => \DATA_OUT_1_15[7]\, DATA_IN_1_15(6)
         => \DATA_OUT_1_15[6]\, DATA_IN_1_15(5) => 
        \DATA_OUT_1_15[5]\, DATA_IN_1_15(4) => \DATA_OUT_1_15[4]\, 
        DATA_IN_1_15(3) => \DATA_OUT_1_15[3]\, DATA_IN_1_15(2)
         => \DATA_OUT_1_15[2]\, DATA_IN_1_15(1) => 
        \DATA_OUT_1_15[1]\, DATA_IN_1_15(0) => \DATA_OUT_1_15[0]\, 
        DATA_IN_1_16(25) => \DATA_OUT_1_16[25]\, DATA_IN_1_16(24)
         => \DATA_OUT_1_16[24]\, DATA_IN_1_16(23) => 
        \DATA_OUT_1_16[23]\, DATA_IN_1_16(22) => 
        \DATA_OUT_1_16[22]\, DATA_IN_1_16(21) => 
        \DATA_OUT_1_16[21]\, DATA_IN_1_16(20) => 
        \DATA_OUT_1_16[20]\, DATA_IN_1_16(19) => 
        \DATA_OUT_1_16[19]\, DATA_IN_1_16(18) => 
        \DATA_OUT_1_16[18]\, DATA_IN_1_16(17) => 
        \DATA_OUT_1_16[17]\, DATA_IN_1_16(16) => 
        \DATA_OUT_1_16[16]\, DATA_IN_1_16(15) => 
        \DATA_OUT_1_16[15]\, DATA_IN_1_16(14) => 
        \DATA_OUT_1_16[14]\, DATA_IN_1_16(13) => 
        \DATA_OUT_1_16[13]\, DATA_IN_1_16(12) => 
        \DATA_OUT_1_16[12]\, DATA_IN_1_16(11) => 
        \DATA_OUT_1_16[11]\, DATA_IN_1_16(10) => 
        \DATA_OUT_1_16[10]\, DATA_IN_1_16(9) => 
        \DATA_OUT_1_16[9]\, DATA_IN_1_16(8) => \DATA_OUT_1_16[8]\, 
        DATA_IN_1_16(7) => \DATA_OUT_1_16[7]\, DATA_IN_1_16(6)
         => \DATA_OUT_1_16[6]\, DATA_IN_1_16(5) => 
        \DATA_OUT_1_16[5]\, DATA_IN_1_16(4) => \DATA_OUT_1_16[4]\, 
        DATA_IN_1_16(3) => \DATA_OUT_1_16[3]\, DATA_IN_1_16(2)
         => \DATA_OUT_1_16[2]\, DATA_IN_1_16(1) => 
        \DATA_OUT_1_16[1]\, DATA_IN_1_16(0) => \DATA_OUT_1_16[0]\, 
        DATA_IN_1_17(25) => \DATA_OUT_1_17[25]\, DATA_IN_1_17(24)
         => \DATA_OUT_1_17[24]\, DATA_IN_1_17(23) => 
        \DATA_OUT_1_17[23]\, DATA_IN_1_17(22) => 
        \DATA_OUT_1_17[22]\, DATA_IN_1_17(21) => 
        \DATA_OUT_1_17[21]\, DATA_IN_1_17(20) => 
        \DATA_OUT_1_17[20]\, DATA_IN_1_17(19) => 
        \DATA_OUT_1_17[19]\, DATA_IN_1_17(18) => 
        \DATA_OUT_1_17[18]\, DATA_IN_1_17(17) => 
        \DATA_OUT_1_17[17]\, DATA_IN_1_17(16) => 
        \DATA_OUT_1_17[16]\, DATA_IN_1_17(15) => 
        \DATA_OUT_1_17[15]\, DATA_IN_1_17(14) => 
        \DATA_OUT_1_17[14]\, DATA_IN_1_17(13) => 
        \DATA_OUT_1_17[13]\, DATA_IN_1_17(12) => 
        \DATA_OUT_1_17[12]\, DATA_IN_1_17(11) => 
        \DATA_OUT_1_17[11]\, DATA_IN_1_17(10) => 
        \DATA_OUT_1_17[10]\, DATA_IN_1_17(9) => 
        \DATA_OUT_1_17[9]\, DATA_IN_1_17(8) => \DATA_OUT_1_17[8]\, 
        DATA_IN_1_17(7) => \DATA_OUT_1_17[7]\, DATA_IN_1_17(6)
         => \DATA_OUT_1_17[6]\, DATA_IN_1_17(5) => 
        \DATA_OUT_1_17[5]\, DATA_IN_1_17(4) => \DATA_OUT_1_17[4]\, 
        DATA_IN_1_17(3) => \DATA_OUT_1_17[3]\, DATA_IN_1_17(2)
         => \DATA_OUT_1_17[2]\, DATA_IN_1_17(1) => 
        \DATA_OUT_1_17[1]\, DATA_IN_1_17(0) => \DATA_OUT_1_17[0]\, 
        DATA_IN_1_18(25) => \DATA_OUT_1_18[25]\, DATA_IN_1_18(24)
         => \DATA_OUT_1_18[24]\, DATA_IN_1_18(23) => 
        \DATA_OUT_1_18[23]\, DATA_IN_1_18(22) => 
        \DATA_OUT_1_18[22]\, DATA_IN_1_18(21) => 
        \DATA_OUT_1_18[21]\, DATA_IN_1_18(20) => 
        \DATA_OUT_1_18[20]\, DATA_IN_1_18(19) => 
        \DATA_OUT_1_18[19]\, DATA_IN_1_18(18) => 
        \DATA_OUT_1_18[18]\, DATA_IN_1_18(17) => 
        \DATA_OUT_1_18[17]\, DATA_IN_1_18(16) => 
        \DATA_OUT_1_18[16]\, DATA_IN_1_18(15) => 
        \DATA_OUT_1_18[15]\, DATA_IN_1_18(14) => 
        \DATA_OUT_1_18[14]\, DATA_IN_1_18(13) => 
        \DATA_OUT_1_18[13]\, DATA_IN_1_18(12) => 
        \DATA_OUT_1_18[12]\, DATA_IN_1_18(11) => 
        \DATA_OUT_1_18[11]\, DATA_IN_1_18(10) => 
        \DATA_OUT_1_18[10]\, DATA_IN_1_18(9) => 
        \DATA_OUT_1_18[9]\, DATA_IN_1_18(8) => \DATA_OUT_1_18[8]\, 
        DATA_IN_1_18(7) => \DATA_OUT_1_18[7]\, DATA_IN_1_18(6)
         => \DATA_OUT_1_18[6]\, DATA_IN_1_18(5) => 
        \DATA_OUT_1_18[5]\, DATA_IN_1_18(4) => \DATA_OUT_1_18[4]\, 
        DATA_IN_1_18(3) => \DATA_OUT_1_18[3]\, DATA_IN_1_18(2)
         => \DATA_OUT_1_18[2]\, DATA_IN_1_18(1) => 
        \DATA_OUT_1_18[1]\, DATA_IN_1_18(0) => \DATA_OUT_1_18[0]\, 
        DATA_IN_1_19(25) => \DATA_OUT_1_19[25]\, DATA_IN_1_19(24)
         => \DATA_OUT_1_19[24]\, DATA_IN_1_19(23) => 
        \DATA_OUT_1_19[23]\, DATA_IN_1_19(22) => 
        \DATA_OUT_1_19[22]\, DATA_IN_1_19(21) => 
        \DATA_OUT_1_19[21]\, DATA_IN_1_19(20) => 
        \DATA_OUT_1_19[20]\, DATA_IN_1_19(19) => 
        \DATA_OUT_1_19[19]\, DATA_IN_1_19(18) => 
        \DATA_OUT_1_19[18]\, DATA_IN_1_19(17) => 
        \DATA_OUT_1_19[17]\, DATA_IN_1_19(16) => 
        \DATA_OUT_1_19[16]\, DATA_IN_1_19(15) => 
        \DATA_OUT_1_19[15]\, DATA_IN_1_19(14) => 
        \DATA_OUT_1_19[14]\, DATA_IN_1_19(13) => 
        \DATA_OUT_1_19[13]\, DATA_IN_1_19(12) => 
        \DATA_OUT_1_19[12]\, DATA_IN_1_19(11) => 
        \DATA_OUT_1_19[11]\, DATA_IN_1_19(10) => 
        \DATA_OUT_1_19[10]\, DATA_IN_1_19(9) => 
        \DATA_OUT_1_19[9]\, DATA_IN_1_19(8) => \DATA_OUT_1_19[8]\, 
        DATA_IN_1_19(7) => \DATA_OUT_1_19[7]\, DATA_IN_1_19(6)
         => \DATA_OUT_1_19[6]\, DATA_IN_1_19(5) => 
        \DATA_OUT_1_19[5]\, DATA_IN_1_19(4) => \DATA_OUT_1_19[4]\, 
        DATA_IN_1_19(3) => \DATA_OUT_1_19[3]\, DATA_IN_1_19(2)
         => \DATA_OUT_1_19[2]\, DATA_IN_1_19(1) => 
        \DATA_OUT_1_19[1]\, DATA_IN_1_19(0) => \DATA_OUT_1_19[0]\, 
        DATA_IN_1_20(25) => \DATA_OUT_1_20[25]\, DATA_IN_1_20(24)
         => \DATA_OUT_1_20[24]\, DATA_IN_1_20(23) => 
        \DATA_OUT_1_20[23]\, DATA_IN_1_20(22) => 
        \DATA_OUT_1_20[22]\, DATA_IN_1_20(21) => 
        \DATA_OUT_1_20[21]\, DATA_IN_1_20(20) => 
        \DATA_OUT_1_20[20]\, DATA_IN_1_20(19) => 
        \DATA_OUT_1_20[19]\, DATA_IN_1_20(18) => 
        \DATA_OUT_1_20[18]\, DATA_IN_1_20(17) => 
        \DATA_OUT_1_20[17]\, DATA_IN_1_20(16) => 
        \DATA_OUT_1_20[16]\, DATA_IN_1_20(15) => 
        \DATA_OUT_1_20[15]\, DATA_IN_1_20(14) => 
        \DATA_OUT_1_20[14]\, DATA_IN_1_20(13) => 
        \DATA_OUT_1_20[13]\, DATA_IN_1_20(12) => 
        \DATA_OUT_1_20[12]\, DATA_IN_1_20(11) => 
        \DATA_OUT_1_20[11]\, DATA_IN_1_20(10) => 
        \DATA_OUT_1_20[10]\, DATA_IN_1_20(9) => 
        \DATA_OUT_1_20[9]\, DATA_IN_1_20(8) => \DATA_OUT_1_20[8]\, 
        DATA_IN_1_20(7) => \DATA_OUT_1_20[7]\, DATA_IN_1_20(6)
         => \DATA_OUT_1_20[6]\, DATA_IN_1_20(5) => 
        \DATA_OUT_1_20[5]\, DATA_IN_1_20(4) => \DATA_OUT_1_20[4]\, 
        DATA_IN_1_20(3) => \DATA_OUT_1_20[3]\, DATA_IN_1_20(2)
         => \DATA_OUT_1_20[2]\, DATA_IN_1_20(1) => 
        \DATA_OUT_1_20[1]\, DATA_IN_1_20(0) => \DATA_OUT_1_20[0]\, 
        DATA_IN_1_21(25) => \DATA_OUT_1_21[25]\, DATA_IN_1_21(24)
         => \DATA_OUT_1_21[24]\, DATA_IN_1_21(23) => 
        \DATA_OUT_1_21[23]\, DATA_IN_1_21(22) => 
        \DATA_OUT_1_21[22]\, DATA_IN_1_21(21) => 
        \DATA_OUT_1_21[21]\, DATA_IN_1_21(20) => 
        \DATA_OUT_1_21[20]\, DATA_IN_1_21(19) => 
        \DATA_OUT_1_21[19]\, DATA_IN_1_21(18) => 
        \DATA_OUT_1_21[18]\, DATA_IN_1_21(17) => 
        \DATA_OUT_1_21[17]\, DATA_IN_1_21(16) => 
        \DATA_OUT_1_21[16]\, DATA_IN_1_21(15) => 
        \DATA_OUT_1_21[15]\, DATA_IN_1_21(14) => 
        \DATA_OUT_1_21[14]\, DATA_IN_1_21(13) => 
        \DATA_OUT_1_21[13]\, DATA_IN_1_21(12) => 
        \DATA_OUT_1_21[12]\, DATA_IN_1_21(11) => 
        \DATA_OUT_1_21[11]\, DATA_IN_1_21(10) => 
        \DATA_OUT_1_21[10]\, DATA_IN_1_21(9) => 
        \DATA_OUT_1_21[9]\, DATA_IN_1_21(8) => \DATA_OUT_1_21[8]\, 
        DATA_IN_1_21(7) => \DATA_OUT_1_21[7]\, DATA_IN_1_21(6)
         => \DATA_OUT_1_21[6]\, DATA_IN_1_21(5) => 
        \DATA_OUT_1_21[5]\, DATA_IN_1_21(4) => \DATA_OUT_1_21[4]\, 
        DATA_IN_1_21(3) => \DATA_OUT_1_21[3]\, DATA_IN_1_21(2)
         => \DATA_OUT_1_21[2]\, DATA_IN_1_21(1) => 
        \DATA_OUT_1_21[1]\, DATA_IN_1_21(0) => \DATA_OUT_1_21[0]\, 
        DATA_IN_1_22(25) => \DATA_OUT_1_22[25]\, DATA_IN_1_22(24)
         => \DATA_OUT_1_22[24]\, DATA_IN_1_22(23) => 
        \DATA_OUT_1_22[23]\, DATA_IN_1_22(22) => 
        \DATA_OUT_1_22[22]\, DATA_IN_1_22(21) => 
        \DATA_OUT_1_22[21]\, DATA_IN_1_22(20) => 
        \DATA_OUT_1_22[20]\, DATA_IN_1_22(19) => 
        \DATA_OUT_1_22[19]\, DATA_IN_1_22(18) => 
        \DATA_OUT_1_22[18]\, DATA_IN_1_22(17) => 
        \DATA_OUT_1_22[17]\, DATA_IN_1_22(16) => 
        \DATA_OUT_1_22[16]\, DATA_IN_1_22(15) => 
        \DATA_OUT_1_22[15]\, DATA_IN_1_22(14) => 
        \DATA_OUT_1_22[14]\, DATA_IN_1_22(13) => 
        \DATA_OUT_1_22[13]\, DATA_IN_1_22(12) => 
        \DATA_OUT_1_22[12]\, DATA_IN_1_22(11) => 
        \DATA_OUT_1_22[11]\, DATA_IN_1_22(10) => 
        \DATA_OUT_1_22[10]\, DATA_IN_1_22(9) => 
        \DATA_OUT_1_22[9]\, DATA_IN_1_22(8) => \DATA_OUT_1_22[8]\, 
        DATA_IN_1_22(7) => \DATA_OUT_1_22[7]\, DATA_IN_1_22(6)
         => \DATA_OUT_1_22[6]\, DATA_IN_1_22(5) => 
        \DATA_OUT_1_22[5]\, DATA_IN_1_22(4) => \DATA_OUT_1_22[4]\, 
        DATA_IN_1_22(3) => \DATA_OUT_1_22[3]\, DATA_IN_1_22(2)
         => \DATA_OUT_1_22[2]\, DATA_IN_1_22(1) => 
        \DATA_OUT_1_22[1]\, DATA_IN_1_22(0) => \DATA_OUT_1_22[0]\, 
        DATA_IN_1_23(25) => \DATA_OUT_1_23[25]\, DATA_IN_1_23(24)
         => \DATA_OUT_1_23[24]\, DATA_IN_1_23(23) => 
        \DATA_OUT_1_23[23]\, DATA_IN_1_23(22) => 
        \DATA_OUT_1_23[22]\, DATA_IN_1_23(21) => 
        \DATA_OUT_1_23[21]\, DATA_IN_1_23(20) => 
        \DATA_OUT_1_23[20]\, DATA_IN_1_23(19) => 
        \DATA_OUT_1_23[19]\, DATA_IN_1_23(18) => 
        \DATA_OUT_1_23[18]\, DATA_IN_1_23(17) => 
        \DATA_OUT_1_23[17]\, DATA_IN_1_23(16) => 
        \DATA_OUT_1_23[16]\, DATA_IN_1_23(15) => 
        \DATA_OUT_1_23[15]\, DATA_IN_1_23(14) => 
        \DATA_OUT_1_23[14]\, DATA_IN_1_23(13) => 
        \DATA_OUT_1_23[13]\, DATA_IN_1_23(12) => 
        \DATA_OUT_1_23[12]\, DATA_IN_1_23(11) => 
        \DATA_OUT_1_23[11]\, DATA_IN_1_23(10) => 
        \DATA_OUT_1_23[10]\, DATA_IN_1_23(9) => 
        \DATA_OUT_1_23[9]\, DATA_IN_1_23(8) => \DATA_OUT_1_23[8]\, 
        DATA_IN_1_23(7) => \DATA_OUT_1_23[7]\, DATA_IN_1_23(6)
         => \DATA_OUT_1_23[6]\, DATA_IN_1_23(5) => 
        \DATA_OUT_1_23[5]\, DATA_IN_1_23(4) => \DATA_OUT_1_23[4]\, 
        DATA_IN_1_23(3) => \DATA_OUT_1_23[3]\, DATA_IN_1_23(2)
         => \DATA_OUT_1_23[2]\, DATA_IN_1_23(1) => 
        \DATA_OUT_1_23[1]\, DATA_IN_1_23(0) => \DATA_OUT_1_23[0]\, 
        DATA_IN_1_24(25) => \DATA_OUT_1_24[25]\, DATA_IN_1_24(24)
         => \DATA_OUT_1_24[24]\, DATA_IN_1_24(23) => 
        \DATA_OUT_1_24[23]\, DATA_IN_1_24(22) => 
        \DATA_OUT_1_24[22]\, DATA_IN_1_24(21) => 
        \DATA_OUT_1_24[21]\, DATA_IN_1_24(20) => 
        \DATA_OUT_1_24[20]\, DATA_IN_1_24(19) => 
        \DATA_OUT_1_24[19]\, DATA_IN_1_24(18) => 
        \DATA_OUT_1_24[18]\, DATA_IN_1_24(17) => 
        \DATA_OUT_1_24[17]\, DATA_IN_1_24(16) => 
        \DATA_OUT_1_24[16]\, DATA_IN_1_24(15) => 
        \DATA_OUT_1_24[15]\, DATA_IN_1_24(14) => 
        \DATA_OUT_1_24[14]\, DATA_IN_1_24(13) => 
        \DATA_OUT_1_24[13]\, DATA_IN_1_24(12) => 
        \DATA_OUT_1_24[12]\, DATA_IN_1_24(11) => 
        \DATA_OUT_1_24[11]\, DATA_IN_1_24(10) => 
        \DATA_OUT_1_24[10]\, DATA_IN_1_24(9) => 
        \DATA_OUT_1_24[9]\, DATA_IN_1_24(8) => \DATA_OUT_1_24[8]\, 
        DATA_IN_1_24(7) => \DATA_OUT_1_24[7]\, DATA_IN_1_24(6)
         => \DATA_OUT_1_24[6]\, DATA_IN_1_24(5) => 
        \DATA_OUT_1_24[5]\, DATA_IN_1_24(4) => \DATA_OUT_1_24[4]\, 
        DATA_IN_1_24(3) => \DATA_OUT_1_24[3]\, DATA_IN_1_24(2)
         => \DATA_OUT_1_24[2]\, DATA_IN_1_24(1) => 
        \DATA_OUT_1_24[1]\, DATA_IN_1_24(0) => \DATA_OUT_1_24[0]\, 
        DATA_IN_1_25(25) => \DATA_OUT_1_25[25]\, DATA_IN_1_25(24)
         => \DATA_OUT_1_25[24]\, DATA_IN_1_25(23) => 
        \DATA_OUT_1_25[23]\, DATA_IN_1_25(22) => 
        \DATA_OUT_1_25[22]\, DATA_IN_1_25(21) => 
        \DATA_OUT_1_25[21]\, DATA_IN_1_25(20) => 
        \DATA_OUT_1_25[20]\, DATA_IN_1_25(19) => 
        \DATA_OUT_1_25[19]\, DATA_IN_1_25(18) => 
        \DATA_OUT_1_25[18]\, DATA_IN_1_25(17) => 
        \DATA_OUT_1_25[17]\, DATA_IN_1_25(16) => 
        \DATA_OUT_1_25[16]\, DATA_IN_1_25(15) => 
        \DATA_OUT_1_25[15]\, DATA_IN_1_25(14) => 
        \DATA_OUT_1_25[14]\, DATA_IN_1_25(13) => 
        \DATA_OUT_1_25[13]\, DATA_IN_1_25(12) => 
        \DATA_OUT_1_25[12]\, DATA_IN_1_25(11) => 
        \DATA_OUT_1_25[11]\, DATA_IN_1_25(10) => 
        \DATA_OUT_1_25[10]\, DATA_IN_1_25(9) => 
        \DATA_OUT_1_25[9]\, DATA_IN_1_25(8) => \DATA_OUT_1_25[8]\, 
        DATA_IN_1_25(7) => \DATA_OUT_1_25[7]\, DATA_IN_1_25(6)
         => \DATA_OUT_1_25[6]\, DATA_IN_1_25(5) => 
        \DATA_OUT_1_25[5]\, DATA_IN_1_25(4) => \DATA_OUT_1_25[4]\, 
        DATA_IN_1_25(3) => \DATA_OUT_1_25[3]\, DATA_IN_1_25(2)
         => \DATA_OUT_1_25[2]\, DATA_IN_1_25(1) => 
        \DATA_OUT_1_25[1]\, DATA_IN_1_25(0) => \DATA_OUT_1_25[0]\, 
        DATA_IN_1_26(25) => \DATA_OUT_1_26[25]\, DATA_IN_1_26(24)
         => \DATA_OUT_1_26[24]\, DATA_IN_1_26(23) => 
        \DATA_OUT_1_26[23]\, DATA_IN_1_26(22) => 
        \DATA_OUT_1_26[22]\, DATA_IN_1_26(21) => 
        \DATA_OUT_1_26[21]\, DATA_IN_1_26(20) => 
        \DATA_OUT_1_26[20]\, DATA_IN_1_26(19) => 
        \DATA_OUT_1_26[19]\, DATA_IN_1_26(18) => 
        \DATA_OUT_1_26[18]\, DATA_IN_1_26(17) => 
        \DATA_OUT_1_26[17]\, DATA_IN_1_26(16) => 
        \DATA_OUT_1_26[16]\, DATA_IN_1_26(15) => 
        \DATA_OUT_1_26[15]\, DATA_IN_1_26(14) => 
        \DATA_OUT_1_26[14]\, DATA_IN_1_26(13) => 
        \DATA_OUT_1_26[13]\, DATA_IN_1_26(12) => 
        \DATA_OUT_1_26[12]\, DATA_IN_1_26(11) => 
        \DATA_OUT_1_26[11]\, DATA_IN_1_26(10) => 
        \DATA_OUT_1_26[10]\, DATA_IN_1_26(9) => 
        \DATA_OUT_1_26[9]\, DATA_IN_1_26(8) => \DATA_OUT_1_26[8]\, 
        DATA_IN_1_26(7) => \DATA_OUT_1_26[7]\, DATA_IN_1_26(6)
         => \DATA_OUT_1_26[6]\, DATA_IN_1_26(5) => 
        \DATA_OUT_1_26[5]\, DATA_IN_1_26(4) => \DATA_OUT_1_26[4]\, 
        DATA_IN_1_26(3) => \DATA_OUT_1_26[3]\, DATA_IN_1_26(2)
         => \DATA_OUT_1_26[2]\, DATA_IN_1_26(1) => 
        \DATA_OUT_1_26[1]\, DATA_IN_1_26(0) => \DATA_OUT_1_26[0]\, 
        DATA_IN_1_27(25) => \DATA_OUT_1_27[25]\, DATA_IN_1_27(24)
         => \DATA_OUT_1_27[24]\, DATA_IN_1_27(23) => 
        \DATA_OUT_1_27[23]\, DATA_IN_1_27(22) => 
        \DATA_OUT_1_27[22]\, DATA_IN_1_27(21) => 
        \DATA_OUT_1_27[21]\, DATA_IN_1_27(20) => 
        \DATA_OUT_1_27[20]\, DATA_IN_1_27(19) => 
        \DATA_OUT_1_27[19]\, DATA_IN_1_27(18) => 
        \DATA_OUT_1_27[18]\, DATA_IN_1_27(17) => 
        \DATA_OUT_1_27[17]\, DATA_IN_1_27(16) => 
        \DATA_OUT_1_27[16]\, DATA_IN_1_27(15) => 
        \DATA_OUT_1_27[15]\, DATA_IN_1_27(14) => 
        \DATA_OUT_1_27[14]\, DATA_IN_1_27(13) => 
        \DATA_OUT_1_27[13]\, DATA_IN_1_27(12) => 
        \DATA_OUT_1_27[12]\, DATA_IN_1_27(11) => 
        \DATA_OUT_1_27[11]\, DATA_IN_1_27(10) => 
        \DATA_OUT_1_27[10]\, DATA_IN_1_27(9) => 
        \DATA_OUT_1_27[9]\, DATA_IN_1_27(8) => \DATA_OUT_1_27[8]\, 
        DATA_IN_1_27(7) => \DATA_OUT_1_27[7]\, DATA_IN_1_27(6)
         => \DATA_OUT_1_27[6]\, DATA_IN_1_27(5) => 
        \DATA_OUT_1_27[5]\, DATA_IN_1_27(4) => \DATA_OUT_1_27[4]\, 
        DATA_IN_1_27(3) => \DATA_OUT_1_27[3]\, DATA_IN_1_27(2)
         => \DATA_OUT_1_27[2]\, DATA_IN_1_27(1) => 
        \DATA_OUT_1_27[1]\, DATA_IN_1_27(0) => \DATA_OUT_1_27[0]\, 
        DATA_IN_1_28(25) => \DATA_OUT_1_28[25]\, DATA_IN_1_28(24)
         => \DATA_OUT_1_28[24]\, DATA_IN_1_28(23) => 
        \DATA_OUT_1_28[23]\, DATA_IN_1_28(22) => 
        \DATA_OUT_1_28[22]\, DATA_IN_1_28(21) => 
        \DATA_OUT_1_28[21]\, DATA_IN_1_28(20) => 
        \DATA_OUT_1_28[20]\, DATA_IN_1_28(19) => 
        \DATA_OUT_1_28[19]\, DATA_IN_1_28(18) => 
        \DATA_OUT_1_28[18]\, DATA_IN_1_28(17) => 
        \DATA_OUT_1_28[17]\, DATA_IN_1_28(16) => 
        \DATA_OUT_1_28[16]\, DATA_IN_1_28(15) => 
        \DATA_OUT_1_28[15]\, DATA_IN_1_28(14) => 
        \DATA_OUT_1_28[14]\, DATA_IN_1_28(13) => 
        \DATA_OUT_1_28[13]\, DATA_IN_1_28(12) => 
        \DATA_OUT_1_28[12]\, DATA_IN_1_28(11) => 
        \DATA_OUT_1_28[11]\, DATA_IN_1_28(10) => 
        \DATA_OUT_1_28[10]\, DATA_IN_1_28(9) => 
        \DATA_OUT_1_28[9]\, DATA_IN_1_28(8) => \DATA_OUT_1_28[8]\, 
        DATA_IN_1_28(7) => \DATA_OUT_1_28[7]\, DATA_IN_1_28(6)
         => \DATA_OUT_1_28[6]\, DATA_IN_1_28(5) => 
        \DATA_OUT_1_28[5]\, DATA_IN_1_28(4) => \DATA_OUT_1_28[4]\, 
        DATA_IN_1_28(3) => \DATA_OUT_1_28[3]\, DATA_IN_1_28(2)
         => \DATA_OUT_1_28[2]\, DATA_IN_1_28(1) => 
        \DATA_OUT_1_28[1]\, DATA_IN_1_28(0) => \DATA_OUT_1_28[0]\, 
        DATA_IN_1_29(25) => \DATA_OUT_1_29[25]\, DATA_IN_1_29(24)
         => \DATA_OUT_1_29[24]\, DATA_IN_1_29(23) => 
        \DATA_OUT_1_29[23]\, DATA_IN_1_29(22) => 
        \DATA_OUT_1_29[22]\, DATA_IN_1_29(21) => 
        \DATA_OUT_1_29[21]\, DATA_IN_1_29(20) => 
        \DATA_OUT_1_29[20]\, DATA_IN_1_29(19) => 
        \DATA_OUT_1_29[19]\, DATA_IN_1_29(18) => 
        \DATA_OUT_1_29[18]\, DATA_IN_1_29(17) => 
        \DATA_OUT_1_29[17]\, DATA_IN_1_29(16) => 
        \DATA_OUT_1_29[16]\, DATA_IN_1_29(15) => 
        \DATA_OUT_1_29[15]\, DATA_IN_1_29(14) => 
        \DATA_OUT_1_29[14]\, DATA_IN_1_29(13) => 
        \DATA_OUT_1_29[13]\, DATA_IN_1_29(12) => 
        \DATA_OUT_1_29[12]\, DATA_IN_1_29(11) => 
        \DATA_OUT_1_29[11]\, DATA_IN_1_29(10) => 
        \DATA_OUT_1_29[10]\, DATA_IN_1_29(9) => 
        \DATA_OUT_1_29[9]\, DATA_IN_1_29(8) => \DATA_OUT_1_29[8]\, 
        DATA_IN_1_29(7) => \DATA_OUT_1_29[7]\, DATA_IN_1_29(6)
         => \DATA_OUT_1_29[6]\, DATA_IN_1_29(5) => 
        \DATA_OUT_1_29[5]\, DATA_IN_1_29(4) => \DATA_OUT_1_29[4]\, 
        DATA_IN_1_29(3) => \DATA_OUT_1_29[3]\, DATA_IN_1_29(2)
         => \DATA_OUT_1_29[2]\, DATA_IN_1_29(1) => 
        \DATA_OUT_1_29[1]\, DATA_IN_1_29(0) => \DATA_OUT_1_29[0]\, 
        DATA_IN_1_30(25) => \DATA_OUT_1_30[25]\, DATA_IN_1_30(24)
         => \DATA_OUT_1_30[24]\, DATA_IN_1_30(23) => 
        \DATA_OUT_1_30[23]\, DATA_IN_1_30(22) => 
        \DATA_OUT_1_30[22]\, DATA_IN_1_30(21) => 
        \DATA_OUT_1_30[21]\, DATA_IN_1_30(20) => 
        \DATA_OUT_1_30[20]\, DATA_IN_1_30(19) => 
        \DATA_OUT_1_30[19]\, DATA_IN_1_30(18) => 
        \DATA_OUT_1_30[18]\, DATA_IN_1_30(17) => 
        \DATA_OUT_1_30[17]\, DATA_IN_1_30(16) => 
        \DATA_OUT_1_30[16]\, DATA_IN_1_30(15) => 
        \DATA_OUT_1_30[15]\, DATA_IN_1_30(14) => 
        \DATA_OUT_1_30[14]\, DATA_IN_1_30(13) => 
        \DATA_OUT_1_30[13]\, DATA_IN_1_30(12) => 
        \DATA_OUT_1_30[12]\, DATA_IN_1_30(11) => 
        \DATA_OUT_1_30[11]\, DATA_IN_1_30(10) => 
        \DATA_OUT_1_30[10]\, DATA_IN_1_30(9) => 
        \DATA_OUT_1_30[9]\, DATA_IN_1_30(8) => \DATA_OUT_1_30[8]\, 
        DATA_IN_1_30(7) => \DATA_OUT_1_30[7]\, DATA_IN_1_30(6)
         => \DATA_OUT_1_30[6]\, DATA_IN_1_30(5) => 
        \DATA_OUT_1_30[5]\, DATA_IN_1_30(4) => \DATA_OUT_1_30[4]\, 
        DATA_IN_1_30(3) => \DATA_OUT_1_30[3]\, DATA_IN_1_30(2)
         => \DATA_OUT_1_30[2]\, DATA_IN_1_30(1) => 
        \DATA_OUT_1_30[1]\, DATA_IN_1_30(0) => \DATA_OUT_1_30[0]\, 
        DATA_IN_1_31(25) => \DATA_OUT_1_31[25]\, DATA_IN_1_31(24)
         => \DATA_OUT_1_31[24]\, DATA_IN_1_31(23) => 
        \DATA_OUT_1_31[23]\, DATA_IN_1_31(22) => 
        \DATA_OUT_1_31[22]\, DATA_IN_1_31(21) => 
        \DATA_OUT_1_31[21]\, DATA_IN_1_31(20) => 
        \DATA_OUT_1_31[20]\, DATA_IN_1_31(19) => 
        \DATA_OUT_1_31[19]\, DATA_IN_1_31(18) => 
        \DATA_OUT_1_31[18]\, DATA_IN_1_31(17) => 
        \DATA_OUT_1_31[17]\, DATA_IN_1_31(16) => 
        \DATA_OUT_1_31[16]\, DATA_IN_1_31(15) => 
        \DATA_OUT_1_31[15]\, DATA_IN_1_31(14) => 
        \DATA_OUT_1_31[14]\, DATA_IN_1_31(13) => 
        \DATA_OUT_1_31[13]\, DATA_IN_1_31(12) => 
        \DATA_OUT_1_31[12]\, DATA_IN_1_31(11) => 
        \DATA_OUT_1_31[11]\, DATA_IN_1_31(10) => 
        \DATA_OUT_1_31[10]\, DATA_IN_1_31(9) => 
        \DATA_OUT_1_31[9]\, DATA_IN_1_31(8) => \DATA_OUT_1_31[8]\, 
        DATA_IN_1_31(7) => \DATA_OUT_1_31[7]\, DATA_IN_1_31(6)
         => \DATA_OUT_1_31[6]\, DATA_IN_1_31(5) => 
        \DATA_OUT_1_31[5]\, DATA_IN_1_31(4) => \DATA_OUT_1_31[4]\, 
        DATA_IN_1_31(3) => \DATA_OUT_1_31[3]\, DATA_IN_1_31(2)
         => \DATA_OUT_1_31[2]\, DATA_IN_1_31(1) => 
        \DATA_OUT_1_31[1]\, DATA_IN_1_31(0) => \DATA_OUT_1_31[0]\, 
        DATA_IN_1_32(25) => \DATA_OUT_1_32[25]\, DATA_IN_1_32(24)
         => \DATA_OUT_1_32[24]\, DATA_IN_1_32(23) => 
        \DATA_OUT_1_32[23]\, DATA_IN_1_32(22) => 
        \DATA_OUT_1_32[22]\, DATA_IN_1_32(21) => 
        \DATA_OUT_1_32[21]\, DATA_IN_1_32(20) => 
        \DATA_OUT_1_32[20]\, DATA_IN_1_32(19) => 
        \DATA_OUT_1_32[19]\, DATA_IN_1_32(18) => 
        \DATA_OUT_1_32[18]\, DATA_IN_1_32(17) => 
        \DATA_OUT_1_32[17]\, DATA_IN_1_32(16) => 
        \DATA_OUT_1_32[16]\, DATA_IN_1_32(15) => 
        \DATA_OUT_1_32[15]\, DATA_IN_1_32(14) => 
        \DATA_OUT_1_32[14]\, DATA_IN_1_32(13) => 
        \DATA_OUT_1_32[13]\, DATA_IN_1_32(12) => 
        \DATA_OUT_1_32[12]\, DATA_IN_1_32(11) => 
        \DATA_OUT_1_32[11]\, DATA_IN_1_32(10) => 
        \DATA_OUT_1_32[10]\, DATA_IN_1_32(9) => 
        \DATA_OUT_1_32[9]\, DATA_IN_1_32(8) => \DATA_OUT_1_32[8]\, 
        DATA_IN_1_32(7) => \DATA_OUT_1_32[7]\, DATA_IN_1_32(6)
         => \DATA_OUT_1_32[6]\, DATA_IN_1_32(5) => 
        \DATA_OUT_1_32[5]\, DATA_IN_1_32(4) => \DATA_OUT_1_32[4]\, 
        DATA_IN_1_32(3) => \DATA_OUT_1_32[3]\, DATA_IN_1_32(2)
         => \DATA_OUT_1_32[2]\, DATA_IN_1_32(1) => 
        \DATA_OUT_1_32[1]\, DATA_IN_1_32(0) => \DATA_OUT_1_32[0]\, 
        DATA_IN_1_33(25) => \DATA_OUT_1_33[25]\, DATA_IN_1_33(24)
         => \DATA_OUT_1_33[24]\, DATA_IN_1_33(23) => 
        \DATA_OUT_1_33[23]\, DATA_IN_1_33(22) => 
        \DATA_OUT_1_33[22]\, DATA_IN_1_33(21) => 
        \DATA_OUT_1_33[21]\, DATA_IN_1_33(20) => 
        \DATA_OUT_1_33[20]\, DATA_IN_1_33(19) => 
        \DATA_OUT_1_33[19]\, DATA_IN_1_33(18) => 
        \DATA_OUT_1_33[18]\, DATA_IN_1_33(17) => 
        \DATA_OUT_1_33[17]\, DATA_IN_1_33(16) => 
        \DATA_OUT_1_33[16]\, DATA_IN_1_33(15) => 
        \DATA_OUT_1_33[15]\, DATA_IN_1_33(14) => 
        \DATA_OUT_1_33[14]\, DATA_IN_1_33(13) => 
        \DATA_OUT_1_33[13]\, DATA_IN_1_33(12) => 
        \DATA_OUT_1_33[12]\, DATA_IN_1_33(11) => 
        \DATA_OUT_1_33[11]\, DATA_IN_1_33(10) => 
        \DATA_OUT_1_33[10]\, DATA_IN_1_33(9) => 
        \DATA_OUT_1_33[9]\, DATA_IN_1_33(8) => \DATA_OUT_1_33[8]\, 
        DATA_IN_1_33(7) => \DATA_OUT_1_33[7]\, DATA_IN_1_33(6)
         => \DATA_OUT_1_33[6]\, DATA_IN_1_33(5) => 
        \DATA_OUT_1_33[5]\, DATA_IN_1_33(4) => \DATA_OUT_1_33[4]\, 
        DATA_IN_1_33(3) => \DATA_OUT_1_33[3]\, DATA_IN_1_33(2)
         => \DATA_OUT_1_33[2]\, DATA_IN_1_33(1) => 
        \DATA_OUT_1_33[1]\, DATA_IN_1_33(0) => \DATA_OUT_1_33[0]\, 
        DATA_IN_1_34(25) => \DATA_OUT_1_34[25]\, DATA_IN_1_34(24)
         => \DATA_OUT_1_34[24]\, DATA_IN_1_34(23) => 
        \DATA_OUT_1_34[23]\, DATA_IN_1_34(22) => 
        \DATA_OUT_1_34[22]\, DATA_IN_1_34(21) => 
        \DATA_OUT_1_34[21]\, DATA_IN_1_34(20) => 
        \DATA_OUT_1_34[20]\, DATA_IN_1_34(19) => 
        \DATA_OUT_1_34[19]\, DATA_IN_1_34(18) => 
        \DATA_OUT_1_34[18]\, DATA_IN_1_34(17) => 
        \DATA_OUT_1_34[17]\, DATA_IN_1_34(16) => 
        \DATA_OUT_1_34[16]\, DATA_IN_1_34(15) => 
        \DATA_OUT_1_34[15]\, DATA_IN_1_34(14) => 
        \DATA_OUT_1_34[14]\, DATA_IN_1_34(13) => 
        \DATA_OUT_1_34[13]\, DATA_IN_1_34(12) => 
        \DATA_OUT_1_34[12]\, DATA_IN_1_34(11) => 
        \DATA_OUT_1_34[11]\, DATA_IN_1_34(10) => 
        \DATA_OUT_1_34[10]\, DATA_IN_1_34(9) => 
        \DATA_OUT_1_34[9]\, DATA_IN_1_34(8) => \DATA_OUT_1_34[8]\, 
        DATA_IN_1_34(7) => \DATA_OUT_1_34[7]\, DATA_IN_1_34(6)
         => \DATA_OUT_1_34[6]\, DATA_IN_1_34(5) => 
        \DATA_OUT_1_34[5]\, DATA_IN_1_34(4) => \DATA_OUT_1_34[4]\, 
        DATA_IN_1_34(3) => \DATA_OUT_1_34[3]\, DATA_IN_1_34(2)
         => \DATA_OUT_1_34[2]\, DATA_IN_1_34(1) => 
        \DATA_OUT_1_34[1]\, DATA_IN_1_34(0) => \DATA_OUT_1_34[0]\, 
        DATA_IN_1_35(25) => \DATA_OUT_1_35[25]\, DATA_IN_1_35(24)
         => \DATA_OUT_1_35[24]\, DATA_IN_1_35(23) => 
        \DATA_OUT_1_35[23]\, DATA_IN_1_35(22) => 
        \DATA_OUT_1_35[22]\, DATA_IN_1_35(21) => 
        \DATA_OUT_1_35[21]\, DATA_IN_1_35(20) => 
        \DATA_OUT_1_35[20]\, DATA_IN_1_35(19) => 
        \DATA_OUT_1_35[19]\, DATA_IN_1_35(18) => 
        \DATA_OUT_1_35[18]\, DATA_IN_1_35(17) => 
        \DATA_OUT_1_35[17]\, DATA_IN_1_35(16) => 
        \DATA_OUT_1_35[16]\, DATA_IN_1_35(15) => 
        \DATA_OUT_1_35[15]\, DATA_IN_1_35(14) => 
        \DATA_OUT_1_35[14]\, DATA_IN_1_35(13) => 
        \DATA_OUT_1_35[13]\, DATA_IN_1_35(12) => 
        \DATA_OUT_1_35[12]\, DATA_IN_1_35(11) => 
        \DATA_OUT_1_35[11]\, DATA_IN_1_35(10) => 
        \DATA_OUT_1_35[10]\, DATA_IN_1_35(9) => 
        \DATA_OUT_1_35[9]\, DATA_IN_1_35(8) => \DATA_OUT_1_35[8]\, 
        DATA_IN_1_35(7) => \DATA_OUT_1_35[7]\, DATA_IN_1_35(6)
         => \DATA_OUT_1_35[6]\, DATA_IN_1_35(5) => 
        \DATA_OUT_1_35[5]\, DATA_IN_1_35(4) => \DATA_OUT_1_35[4]\, 
        DATA_IN_1_35(3) => \DATA_OUT_1_35[3]\, DATA_IN_1_35(2)
         => \DATA_OUT_1_35[2]\, DATA_IN_1_35(1) => 
        \DATA_OUT_1_35[1]\, DATA_IN_1_35(0) => \DATA_OUT_1_35[0]\, 
        DATA_IN_1_36(25) => \DATA_OUT_1_36[25]\, DATA_IN_1_36(24)
         => \DATA_OUT_1_36[24]\, DATA_IN_1_36(23) => 
        \DATA_OUT_1_36[23]\, DATA_IN_1_36(22) => 
        \DATA_OUT_1_36[22]\, DATA_IN_1_36(21) => 
        \DATA_OUT_1_36[21]\, DATA_IN_1_36(20) => 
        \DATA_OUT_1_36[20]\, DATA_IN_1_36(19) => 
        \DATA_OUT_1_36[19]\, DATA_IN_1_36(18) => 
        \DATA_OUT_1_36[18]\, DATA_IN_1_36(17) => 
        \DATA_OUT_1_36[17]\, DATA_IN_1_36(16) => 
        \DATA_OUT_1_36[16]\, DATA_IN_1_36(15) => 
        \DATA_OUT_1_36[15]\, DATA_IN_1_36(14) => 
        \DATA_OUT_1_36[14]\, DATA_IN_1_36(13) => 
        \DATA_OUT_1_36[13]\, DATA_IN_1_36(12) => 
        \DATA_OUT_1_36[12]\, DATA_IN_1_36(11) => 
        \DATA_OUT_1_36[11]\, DATA_IN_1_36(10) => 
        \DATA_OUT_1_36[10]\, DATA_IN_1_36(9) => 
        \DATA_OUT_1_36[9]\, DATA_IN_1_36(8) => \DATA_OUT_1_36[8]\, 
        DATA_IN_1_36(7) => \DATA_OUT_1_36[7]\, DATA_IN_1_36(6)
         => \DATA_OUT_1_36[6]\, DATA_IN_1_36(5) => 
        \DATA_OUT_1_36[5]\, DATA_IN_1_36(4) => \DATA_OUT_1_36[4]\, 
        DATA_IN_1_36(3) => \DATA_OUT_1_36[3]\, DATA_IN_1_36(2)
         => \DATA_OUT_1_36[2]\, DATA_IN_1_36(1) => 
        \DATA_OUT_1_36[1]\, DATA_IN_1_36(0) => \DATA_OUT_1_36[0]\, 
        DATA_IN_1_37(25) => \DATA_OUT_1_37[25]\, DATA_IN_1_37(24)
         => \DATA_OUT_1_37[24]\, DATA_IN_1_37(23) => 
        \DATA_OUT_1_37[23]\, DATA_IN_1_37(22) => 
        \DATA_OUT_1_37[22]\, DATA_IN_1_37(21) => 
        \DATA_OUT_1_37[21]\, DATA_IN_1_37(20) => 
        \DATA_OUT_1_37[20]\, DATA_IN_1_37(19) => 
        \DATA_OUT_1_37[19]\, DATA_IN_1_37(18) => 
        \DATA_OUT_1_37[18]\, DATA_IN_1_37(17) => 
        \DATA_OUT_1_37[17]\, DATA_IN_1_37(16) => 
        \DATA_OUT_1_37[16]\, DATA_IN_1_37(15) => 
        \DATA_OUT_1_37[15]\, DATA_IN_1_37(14) => 
        \DATA_OUT_1_37[14]\, DATA_IN_1_37(13) => 
        \DATA_OUT_1_37[13]\, DATA_IN_1_37(12) => 
        \DATA_OUT_1_37[12]\, DATA_IN_1_37(11) => 
        \DATA_OUT_1_37[11]\, DATA_IN_1_37(10) => 
        \DATA_OUT_1_37[10]\, DATA_IN_1_37(9) => 
        \DATA_OUT_1_37[9]\, DATA_IN_1_37(8) => \DATA_OUT_1_37[8]\, 
        DATA_IN_1_37(7) => \DATA_OUT_1_37[7]\, DATA_IN_1_37(6)
         => \DATA_OUT_1_37[6]\, DATA_IN_1_37(5) => 
        \DATA_OUT_1_37[5]\, DATA_IN_1_37(4) => \DATA_OUT_1_37[4]\, 
        DATA_IN_1_37(3) => \DATA_OUT_1_37[3]\, DATA_IN_1_37(2)
         => \DATA_OUT_1_37[2]\, DATA_IN_1_37(1) => 
        \DATA_OUT_1_37[1]\, DATA_IN_1_37(0) => \DATA_OUT_1_37[0]\, 
        DATA_IN_1_38(25) => \DATA_OUT_1_38[25]\, DATA_IN_1_38(24)
         => \DATA_OUT_1_38[24]\, DATA_IN_1_38(23) => 
        \DATA_OUT_1_38[23]\, DATA_IN_1_38(22) => 
        \DATA_OUT_1_38[22]\, DATA_IN_1_38(21) => 
        \DATA_OUT_1_38[21]\, DATA_IN_1_38(20) => 
        \DATA_OUT_1_38[20]\, DATA_IN_1_38(19) => 
        \DATA_OUT_1_38[19]\, DATA_IN_1_38(18) => 
        \DATA_OUT_1_38[18]\, DATA_IN_1_38(17) => 
        \DATA_OUT_1_38[17]\, DATA_IN_1_38(16) => 
        \DATA_OUT_1_38[16]\, DATA_IN_1_38(15) => 
        \DATA_OUT_1_38[15]\, DATA_IN_1_38(14) => 
        \DATA_OUT_1_38[14]\, DATA_IN_1_38(13) => 
        \DATA_OUT_1_38[13]\, DATA_IN_1_38(12) => 
        \DATA_OUT_1_38[12]\, DATA_IN_1_38(11) => 
        \DATA_OUT_1_38[11]\, DATA_IN_1_38(10) => 
        \DATA_OUT_1_38[10]\, DATA_IN_1_38(9) => 
        \DATA_OUT_1_38[9]\, DATA_IN_1_38(8) => \DATA_OUT_1_38[8]\, 
        DATA_IN_1_38(7) => \DATA_OUT_1_38[7]\, DATA_IN_1_38(6)
         => \DATA_OUT_1_38[6]\, DATA_IN_1_38(5) => 
        \DATA_OUT_1_38[5]\, DATA_IN_1_38(4) => \DATA_OUT_1_38[4]\, 
        DATA_IN_1_38(3) => \DATA_OUT_1_38[3]\, DATA_IN_1_38(2)
         => \DATA_OUT_1_38[2]\, DATA_IN_1_38(1) => 
        \DATA_OUT_1_38[1]\, DATA_IN_1_38(0) => \DATA_OUT_1_38[0]\, 
        DATA_IN_1_39(25) => \DATA_OUT_1_39[25]\, DATA_IN_1_39(24)
         => \DATA_OUT_1_39[24]\, DATA_IN_1_39(23) => 
        \DATA_OUT_1_39[23]\, DATA_IN_1_39(22) => 
        \DATA_OUT_1_39[22]\, DATA_IN_1_39(21) => 
        \DATA_OUT_1_39[21]\, DATA_IN_1_39(20) => 
        \DATA_OUT_1_39[20]\, DATA_IN_1_39(19) => 
        \DATA_OUT_1_39[19]\, DATA_IN_1_39(18) => 
        \DATA_OUT_1_39[18]\, DATA_IN_1_39(17) => 
        \DATA_OUT_1_39[17]\, DATA_IN_1_39(16) => 
        \DATA_OUT_1_39[16]\, DATA_IN_1_39(15) => 
        \DATA_OUT_1_39[15]\, DATA_IN_1_39(14) => 
        \DATA_OUT_1_39[14]\, DATA_IN_1_39(13) => 
        \DATA_OUT_1_39[13]\, DATA_IN_1_39(12) => 
        \DATA_OUT_1_39[12]\, DATA_IN_1_39(11) => 
        \DATA_OUT_1_39[11]\, DATA_IN_1_39(10) => 
        \DATA_OUT_1_39[10]\, DATA_IN_1_39(9) => 
        \DATA_OUT_1_39[9]\, DATA_IN_1_39(8) => \DATA_OUT_1_39[8]\, 
        DATA_IN_1_39(7) => \DATA_OUT_1_39[7]\, DATA_IN_1_39(6)
         => \DATA_OUT_1_39[6]\, DATA_IN_1_39(5) => 
        \DATA_OUT_1_39[5]\, DATA_IN_1_39(4) => \DATA_OUT_1_39[4]\, 
        DATA_IN_1_39(3) => \DATA_OUT_1_39[3]\, DATA_IN_1_39(2)
         => \DATA_OUT_1_39[2]\, DATA_IN_1_39(1) => 
        \DATA_OUT_1_39[1]\, DATA_IN_1_39(0) => \DATA_OUT_1_39[0]\, 
        DATA_IN_1_40(25) => \DATA_OUT_1_40[25]\, DATA_IN_1_40(24)
         => \DATA_OUT_1_40[24]\, DATA_IN_1_40(23) => 
        \DATA_OUT_1_40[23]\, DATA_IN_1_40(22) => 
        \DATA_OUT_1_40[22]\, DATA_IN_1_40(21) => 
        \DATA_OUT_1_40[21]\, DATA_IN_1_40(20) => 
        \DATA_OUT_1_40[20]\, DATA_IN_1_40(19) => 
        \DATA_OUT_1_40[19]\, DATA_IN_1_40(18) => 
        \DATA_OUT_1_40[18]\, DATA_IN_1_40(17) => 
        \DATA_OUT_1_40[17]\, DATA_IN_1_40(16) => 
        \DATA_OUT_1_40[16]\, DATA_IN_1_40(15) => 
        \DATA_OUT_1_40[15]\, DATA_IN_1_40(14) => 
        \DATA_OUT_1_40[14]\, DATA_IN_1_40(13) => 
        \DATA_OUT_1_40[13]\, DATA_IN_1_40(12) => 
        \DATA_OUT_1_40[12]\, DATA_IN_1_40(11) => 
        \DATA_OUT_1_40[11]\, DATA_IN_1_40(10) => 
        \DATA_OUT_1_40[10]\, DATA_IN_1_40(9) => 
        \DATA_OUT_1_40[9]\, DATA_IN_1_40(8) => \DATA_OUT_1_40[8]\, 
        DATA_IN_1_40(7) => \DATA_OUT_1_40[7]\, DATA_IN_1_40(6)
         => \DATA_OUT_1_40[6]\, DATA_IN_1_40(5) => 
        \DATA_OUT_1_40[5]\, DATA_IN_1_40(4) => \DATA_OUT_1_40[4]\, 
        DATA_IN_1_40(3) => \DATA_OUT_1_40[3]\, DATA_IN_1_40(2)
         => \DATA_OUT_1_40[2]\, DATA_IN_1_40(1) => 
        \DATA_OUT_1_40[1]\, DATA_IN_1_40(0) => \DATA_OUT_1_40[0]\, 
        DATA_IN_1_41(25) => \DATA_OUT_1_41[25]\, DATA_IN_1_41(24)
         => \DATA_OUT_1_41[24]\, DATA_IN_1_41(23) => 
        \DATA_OUT_1_41[23]\, DATA_IN_1_41(22) => 
        \DATA_OUT_1_41[22]\, DATA_IN_1_41(21) => 
        \DATA_OUT_1_41[21]\, DATA_IN_1_41(20) => 
        \DATA_OUT_1_41[20]\, DATA_IN_1_41(19) => 
        \DATA_OUT_1_41[19]\, DATA_IN_1_41(18) => 
        \DATA_OUT_1_41[18]\, DATA_IN_1_41(17) => 
        \DATA_OUT_1_41[17]\, DATA_IN_1_41(16) => 
        \DATA_OUT_1_41[16]\, DATA_IN_1_41(15) => 
        \DATA_OUT_1_41[15]\, DATA_IN_1_41(14) => 
        \DATA_OUT_1_41[14]\, DATA_IN_1_41(13) => 
        \DATA_OUT_1_41[13]\, DATA_IN_1_41(12) => 
        \DATA_OUT_1_41[12]\, DATA_IN_1_41(11) => 
        \DATA_OUT_1_41[11]\, DATA_IN_1_41(10) => 
        \DATA_OUT_1_41[10]\, DATA_IN_1_41(9) => 
        \DATA_OUT_1_41[9]\, DATA_IN_1_41(8) => \DATA_OUT_1_41[8]\, 
        DATA_IN_1_41(7) => \DATA_OUT_1_41[7]\, DATA_IN_1_41(6)
         => \DATA_OUT_1_41[6]\, DATA_IN_1_41(5) => 
        \DATA_OUT_1_41[5]\, DATA_IN_1_41(4) => \DATA_OUT_1_41[4]\, 
        DATA_IN_1_41(3) => \DATA_OUT_1_41[3]\, DATA_IN_1_41(2)
         => \DATA_OUT_1_41[2]\, DATA_IN_1_41(1) => 
        \DATA_OUT_1_41[1]\, DATA_IN_1_41(0) => \DATA_OUT_1_41[0]\, 
        DATA_IN_1_42(25) => \DATA_OUT_1_42[25]\, DATA_IN_1_42(24)
         => \DATA_OUT_1_42[24]\, DATA_IN_1_42(23) => 
        \DATA_OUT_1_42[23]\, DATA_IN_1_42(22) => 
        \DATA_OUT_1_42[22]\, DATA_IN_1_42(21) => 
        \DATA_OUT_1_42[21]\, DATA_IN_1_42(20) => 
        \DATA_OUT_1_42[20]\, DATA_IN_1_42(19) => 
        \DATA_OUT_1_42[19]\, DATA_IN_1_42(18) => 
        \DATA_OUT_1_42[18]\, DATA_IN_1_42(17) => 
        \DATA_OUT_1_42[17]\, DATA_IN_1_42(16) => 
        \DATA_OUT_1_42[16]\, DATA_IN_1_42(15) => 
        \DATA_OUT_1_42[15]\, DATA_IN_1_42(14) => 
        \DATA_OUT_1_42[14]\, DATA_IN_1_42(13) => 
        \DATA_OUT_1_42[13]\, DATA_IN_1_42(12) => 
        \DATA_OUT_1_42[12]\, DATA_IN_1_42(11) => 
        \DATA_OUT_1_42[11]\, DATA_IN_1_42(10) => 
        \DATA_OUT_1_42[10]\, DATA_IN_1_42(9) => 
        \DATA_OUT_1_42[9]\, DATA_IN_1_42(8) => \DATA_OUT_1_42[8]\, 
        DATA_IN_1_42(7) => \DATA_OUT_1_42[7]\, DATA_IN_1_42(6)
         => \DATA_OUT_1_42[6]\, DATA_IN_1_42(5) => 
        \DATA_OUT_1_42[5]\, DATA_IN_1_42(4) => \DATA_OUT_1_42[4]\, 
        DATA_IN_1_42(3) => \DATA_OUT_1_42[3]\, DATA_IN_1_42(2)
         => \DATA_OUT_1_42[2]\, DATA_IN_1_42(1) => 
        \DATA_OUT_1_42[1]\, DATA_IN_1_42(0) => \DATA_OUT_1_42[0]\, 
        DATA_IN_1_43(25) => \DATA_OUT_1_43[25]\, DATA_IN_1_43(24)
         => \DATA_OUT_1_43[24]\, DATA_IN_1_43(23) => 
        \DATA_OUT_1_43[23]\, DATA_IN_1_43(22) => 
        \DATA_OUT_1_43[22]\, DATA_IN_1_43(21) => 
        \DATA_OUT_1_43[21]\, DATA_IN_1_43(20) => 
        \DATA_OUT_1_43[20]\, DATA_IN_1_43(19) => 
        \DATA_OUT_1_43[19]\, DATA_IN_1_43(18) => 
        \DATA_OUT_1_43[18]\, DATA_IN_1_43(17) => 
        \DATA_OUT_1_43[17]\, DATA_IN_1_43(16) => 
        \DATA_OUT_1_43[16]\, DATA_IN_1_43(15) => 
        \DATA_OUT_1_43[15]\, DATA_IN_1_43(14) => 
        \DATA_OUT_1_43[14]\, DATA_IN_1_43(13) => 
        \DATA_OUT_1_43[13]\, DATA_IN_1_43(12) => 
        \DATA_OUT_1_43[12]\, DATA_IN_1_43(11) => 
        \DATA_OUT_1_43[11]\, DATA_IN_1_43(10) => 
        \DATA_OUT_1_43[10]\, DATA_IN_1_43(9) => 
        \DATA_OUT_1_43[9]\, DATA_IN_1_43(8) => \DATA_OUT_1_43[8]\, 
        DATA_IN_1_43(7) => \DATA_OUT_1_43[7]\, DATA_IN_1_43(6)
         => \DATA_OUT_1_43[6]\, DATA_IN_1_43(5) => 
        \DATA_OUT_1_43[5]\, DATA_IN_1_43(4) => \DATA_OUT_1_43[4]\, 
        DATA_IN_1_43(3) => \DATA_OUT_1_43[3]\, DATA_IN_1_43(2)
         => \DATA_OUT_1_43[2]\, DATA_IN_1_43(1) => 
        \DATA_OUT_1_43[1]\, DATA_IN_1_43(0) => \DATA_OUT_1_43[0]\, 
        DATA_IN_1_44(25) => \DATA_OUT_1_44[25]\, DATA_IN_1_44(24)
         => \DATA_OUT_1_44[24]\, DATA_IN_1_44(23) => 
        \DATA_OUT_1_44[23]\, DATA_IN_1_44(22) => 
        \DATA_OUT_1_44[22]\, DATA_IN_1_44(21) => 
        \DATA_OUT_1_44[21]\, DATA_IN_1_44(20) => 
        \DATA_OUT_1_44[20]\, DATA_IN_1_44(19) => 
        \DATA_OUT_1_44[19]\, DATA_IN_1_44(18) => 
        \DATA_OUT_1_44[18]\, DATA_IN_1_44(17) => 
        \DATA_OUT_1_44[17]\, DATA_IN_1_44(16) => 
        \DATA_OUT_1_44[16]\, DATA_IN_1_44(15) => 
        \DATA_OUT_1_44[15]\, DATA_IN_1_44(14) => 
        \DATA_OUT_1_44[14]\, DATA_IN_1_44(13) => 
        \DATA_OUT_1_44[13]\, DATA_IN_1_44(12) => 
        \DATA_OUT_1_44[12]\, DATA_IN_1_44(11) => 
        \DATA_OUT_1_44[11]\, DATA_IN_1_44(10) => 
        \DATA_OUT_1_44[10]\, DATA_IN_1_44(9) => 
        \DATA_OUT_1_44[9]\, DATA_IN_1_44(8) => \DATA_OUT_1_44[8]\, 
        DATA_IN_1_44(7) => \DATA_OUT_1_44[7]\, DATA_IN_1_44(6)
         => \DATA_OUT_1_44[6]\, DATA_IN_1_44(5) => 
        \DATA_OUT_1_44[5]\, DATA_IN_1_44(4) => \DATA_OUT_1_44[4]\, 
        DATA_IN_1_44(3) => \DATA_OUT_1_44[3]\, DATA_IN_1_44(2)
         => \DATA_OUT_1_44[2]\, DATA_IN_1_44(1) => 
        \DATA_OUT_1_44[1]\, DATA_IN_1_44(0) => \DATA_OUT_1_44[0]\, 
        DATA_IN_1_45(25) => \DATA_OUT_1_45[25]\, DATA_IN_1_45(24)
         => \DATA_OUT_1_45[24]\, DATA_IN_1_45(23) => 
        \DATA_OUT_1_45[23]\, DATA_IN_1_45(22) => 
        \DATA_OUT_1_45[22]\, DATA_IN_1_45(21) => 
        \DATA_OUT_1_45[21]\, DATA_IN_1_45(20) => 
        \DATA_OUT_1_45[20]\, DATA_IN_1_45(19) => 
        \DATA_OUT_1_45[19]\, DATA_IN_1_45(18) => 
        \DATA_OUT_1_45[18]\, DATA_IN_1_45(17) => 
        \DATA_OUT_1_45[17]\, DATA_IN_1_45(16) => 
        \DATA_OUT_1_45[16]\, DATA_IN_1_45(15) => 
        \DATA_OUT_1_45[15]\, DATA_IN_1_45(14) => 
        \DATA_OUT_1_45[14]\, DATA_IN_1_45(13) => 
        \DATA_OUT_1_45[13]\, DATA_IN_1_45(12) => 
        \DATA_OUT_1_45[12]\, DATA_IN_1_45(11) => 
        \DATA_OUT_1_45[11]\, DATA_IN_1_45(10) => 
        \DATA_OUT_1_45[10]\, DATA_IN_1_45(9) => 
        \DATA_OUT_1_45[9]\, DATA_IN_1_45(8) => \DATA_OUT_1_45[8]\, 
        DATA_IN_1_45(7) => \DATA_OUT_1_45[7]\, DATA_IN_1_45(6)
         => \DATA_OUT_1_45[6]\, DATA_IN_1_45(5) => 
        \DATA_OUT_1_45[5]\, DATA_IN_1_45(4) => \DATA_OUT_1_45[4]\, 
        DATA_IN_1_45(3) => \DATA_OUT_1_45[3]\, DATA_IN_1_45(2)
         => \DATA_OUT_1_45[2]\, DATA_IN_1_45(1) => 
        \DATA_OUT_1_45[1]\, DATA_IN_1_45(0) => \DATA_OUT_1_45[0]\, 
        DATA_IN_1_46(25) => \DATA_OUT_1_46[25]\, DATA_IN_1_46(24)
         => \DATA_OUT_1_46[24]\, DATA_IN_1_46(23) => 
        \DATA_OUT_1_46[23]\, DATA_IN_1_46(22) => 
        \DATA_OUT_1_46[22]\, DATA_IN_1_46(21) => 
        \DATA_OUT_1_46[21]\, DATA_IN_1_46(20) => 
        \DATA_OUT_1_46[20]\, DATA_IN_1_46(19) => 
        \DATA_OUT_1_46[19]\, DATA_IN_1_46(18) => 
        \DATA_OUT_1_46[18]\, DATA_IN_1_46(17) => 
        \DATA_OUT_1_46[17]\, DATA_IN_1_46(16) => 
        \DATA_OUT_1_46[16]\, DATA_IN_1_46(15) => 
        \DATA_OUT_1_46[15]\, DATA_IN_1_46(14) => 
        \DATA_OUT_1_46[14]\, DATA_IN_1_46(13) => 
        \DATA_OUT_1_46[13]\, DATA_IN_1_46(12) => 
        \DATA_OUT_1_46[12]\, DATA_IN_1_46(11) => 
        \DATA_OUT_1_46[11]\, DATA_IN_1_46(10) => 
        \DATA_OUT_1_46[10]\, DATA_IN_1_46(9) => 
        \DATA_OUT_1_46[9]\, DATA_IN_1_46(8) => \DATA_OUT_1_46[8]\, 
        DATA_IN_1_46(7) => \DATA_OUT_1_46[7]\, DATA_IN_1_46(6)
         => \DATA_OUT_1_46[6]\, DATA_IN_1_46(5) => 
        \DATA_OUT_1_46[5]\, DATA_IN_1_46(4) => \DATA_OUT_1_46[4]\, 
        DATA_IN_1_46(3) => \DATA_OUT_1_46[3]\, DATA_IN_1_46(2)
         => \DATA_OUT_1_46[2]\, DATA_IN_1_46(1) => 
        \DATA_OUT_1_46[1]\, DATA_IN_1_46(0) => \DATA_OUT_1_46[0]\, 
        DATA_IN_1_47(25) => \DATA_OUT_1_47[25]\, DATA_IN_1_47(24)
         => \DATA_OUT_1_47[24]\, DATA_IN_1_47(23) => 
        \DATA_OUT_1_47[23]\, DATA_IN_1_47(22) => 
        \DATA_OUT_1_47[22]\, DATA_IN_1_47(21) => 
        \DATA_OUT_1_47[21]\, DATA_IN_1_47(20) => 
        \DATA_OUT_1_47[20]\, DATA_IN_1_47(19) => 
        \DATA_OUT_1_47[19]\, DATA_IN_1_47(18) => 
        \DATA_OUT_1_47[18]\, DATA_IN_1_47(17) => 
        \DATA_OUT_1_47[17]\, DATA_IN_1_47(16) => 
        \DATA_OUT_1_47[16]\, DATA_IN_1_47(15) => 
        \DATA_OUT_1_47[15]\, DATA_IN_1_47(14) => 
        \DATA_OUT_1_47[14]\, DATA_IN_1_47(13) => 
        \DATA_OUT_1_47[13]\, DATA_IN_1_47(12) => 
        \DATA_OUT_1_47[12]\, DATA_IN_1_47(11) => 
        \DATA_OUT_1_47[11]\, DATA_IN_1_47(10) => 
        \DATA_OUT_1_47[10]\, DATA_IN_1_47(9) => 
        \DATA_OUT_1_47[9]\, DATA_IN_1_47(8) => \DATA_OUT_1_47[8]\, 
        DATA_IN_1_47(7) => \DATA_OUT_1_47[7]\, DATA_IN_1_47(6)
         => \DATA_OUT_1_47[6]\, DATA_IN_1_47(5) => 
        \DATA_OUT_1_47[5]\, DATA_IN_1_47(4) => \DATA_OUT_1_47[4]\, 
        DATA_IN_1_47(3) => \DATA_OUT_1_47[3]\, DATA_IN_1_47(2)
         => \DATA_OUT_1_47[2]\, DATA_IN_1_47(1) => 
        \DATA_OUT_1_47[1]\, DATA_IN_1_47(0) => \DATA_OUT_1_47[0]\, 
        DATA_IN_1_48(25) => \DATA_OUT_1_48[25]\, DATA_IN_1_48(24)
         => \DATA_OUT_1_48[24]\, DATA_IN_1_48(23) => 
        \DATA_OUT_1_48[23]\, DATA_IN_1_48(22) => 
        \DATA_OUT_1_48[22]\, DATA_IN_1_48(21) => 
        \DATA_OUT_1_48[21]\, DATA_IN_1_48(20) => 
        \DATA_OUT_1_48[20]\, DATA_IN_1_48(19) => 
        \DATA_OUT_1_48[19]\, DATA_IN_1_48(18) => 
        \DATA_OUT_1_48[18]\, DATA_IN_1_48(17) => 
        \DATA_OUT_1_48[17]\, DATA_IN_1_48(16) => 
        \DATA_OUT_1_48[16]\, DATA_IN_1_48(15) => 
        \DATA_OUT_1_48[15]\, DATA_IN_1_48(14) => 
        \DATA_OUT_1_48[14]\, DATA_IN_1_48(13) => 
        \DATA_OUT_1_48[13]\, DATA_IN_1_48(12) => 
        \DATA_OUT_1_48[12]\, DATA_IN_1_48(11) => 
        \DATA_OUT_1_48[11]\, DATA_IN_1_48(10) => 
        \DATA_OUT_1_48[10]\, DATA_IN_1_48(9) => 
        \DATA_OUT_1_48[9]\, DATA_IN_1_48(8) => \DATA_OUT_1_48[8]\, 
        DATA_IN_1_48(7) => \DATA_OUT_1_48[7]\, DATA_IN_1_48(6)
         => \DATA_OUT_1_48[6]\, DATA_IN_1_48(5) => 
        \DATA_OUT_1_48[5]\, DATA_IN_1_48(4) => \DATA_OUT_1_48[4]\, 
        DATA_IN_1_48(3) => \DATA_OUT_1_48[3]\, DATA_IN_1_48(2)
         => \DATA_OUT_1_48[2]\, DATA_IN_1_48(1) => 
        \DATA_OUT_1_48[1]\, DATA_IN_1_48(0) => \DATA_OUT_1_48[0]\, 
        DATA_IN_1_49(25) => \DATA_OUT_1_49[25]\, DATA_IN_1_49(24)
         => \DATA_OUT_1_49[24]\, DATA_IN_1_49(23) => 
        \DATA_OUT_1_49[23]\, DATA_IN_1_49(22) => 
        \DATA_OUT_1_49[22]\, DATA_IN_1_49(21) => 
        \DATA_OUT_1_49[21]\, DATA_IN_1_49(20) => 
        \DATA_OUT_1_49[20]\, DATA_IN_1_49(19) => 
        \DATA_OUT_1_49[19]\, DATA_IN_1_49(18) => 
        \DATA_OUT_1_49[18]\, DATA_IN_1_49(17) => 
        \DATA_OUT_1_49[17]\, DATA_IN_1_49(16) => 
        \DATA_OUT_1_49[16]\, DATA_IN_1_49(15) => 
        \DATA_OUT_1_49[15]\, DATA_IN_1_49(14) => 
        \DATA_OUT_1_49[14]\, DATA_IN_1_49(13) => 
        \DATA_OUT_1_49[13]\, DATA_IN_1_49(12) => 
        \DATA_OUT_1_49[12]\, DATA_IN_1_49(11) => 
        \DATA_OUT_1_49[11]\, DATA_IN_1_49(10) => 
        \DATA_OUT_1_49[10]\, DATA_IN_1_49(9) => 
        \DATA_OUT_1_49[9]\, DATA_IN_1_49(8) => \DATA_OUT_1_49[8]\, 
        DATA_IN_1_49(7) => \DATA_OUT_1_49[7]\, DATA_IN_1_49(6)
         => \DATA_OUT_1_49[6]\, DATA_IN_1_49(5) => 
        \DATA_OUT_1_49[5]\, DATA_IN_1_49(4) => \DATA_OUT_1_49[4]\, 
        DATA_IN_1_49(3) => \DATA_OUT_1_49[3]\, DATA_IN_1_49(2)
         => \DATA_OUT_1_49[2]\, DATA_IN_1_49(1) => 
        \DATA_OUT_1_49[1]\, DATA_IN_1_49(0) => \DATA_OUT_1_49[0]\, 
        DATA_IN_1_50(25) => \DATA_OUT_1_50[25]\, DATA_IN_1_50(24)
         => \DATA_OUT_1_50[24]\, DATA_IN_1_50(23) => 
        \DATA_OUT_1_50[23]\, DATA_IN_1_50(22) => 
        \DATA_OUT_1_50[22]\, DATA_IN_1_50(21) => 
        \DATA_OUT_1_50[21]\, DATA_IN_1_50(20) => 
        \DATA_OUT_1_50[20]\, DATA_IN_1_50(19) => 
        \DATA_OUT_1_50[19]\, DATA_IN_1_50(18) => 
        \DATA_OUT_1_50[18]\, DATA_IN_1_50(17) => 
        \DATA_OUT_1_50[17]\, DATA_IN_1_50(16) => 
        \DATA_OUT_1_50[16]\, DATA_IN_1_50(15) => 
        \DATA_OUT_1_50[15]\, DATA_IN_1_50(14) => 
        \DATA_OUT_1_50[14]\, DATA_IN_1_50(13) => 
        \DATA_OUT_1_50[13]\, DATA_IN_1_50(12) => 
        \DATA_OUT_1_50[12]\, DATA_IN_1_50(11) => 
        \DATA_OUT_1_50[11]\, DATA_IN_1_50(10) => 
        \DATA_OUT_1_50[10]\, DATA_IN_1_50(9) => 
        \DATA_OUT_1_50[9]\, DATA_IN_1_50(8) => \DATA_OUT_1_50[8]\, 
        DATA_IN_1_50(7) => \DATA_OUT_1_50[7]\, DATA_IN_1_50(6)
         => \DATA_OUT_1_50[6]\, DATA_IN_1_50(5) => 
        \DATA_OUT_1_50[5]\, DATA_IN_1_50(4) => \DATA_OUT_1_50[4]\, 
        DATA_IN_1_50(3) => \DATA_OUT_1_50[3]\, DATA_IN_1_50(2)
         => \DATA_OUT_1_50[2]\, DATA_IN_1_50(1) => 
        \DATA_OUT_1_50[1]\, DATA_IN_1_50(0) => \DATA_OUT_1_50[0]\, 
        DATA_IN_1_51(25) => \DATA_OUT_1_51[25]\, DATA_IN_1_51(24)
         => \DATA_OUT_1_51[24]\, DATA_IN_1_51(23) => 
        \DATA_OUT_1_51[23]\, DATA_IN_1_51(22) => 
        \DATA_OUT_1_51[22]\, DATA_IN_1_51(21) => 
        \DATA_OUT_1_51[21]\, DATA_IN_1_51(20) => 
        \DATA_OUT_1_51[20]\, DATA_IN_1_51(19) => 
        \DATA_OUT_1_51[19]\, DATA_IN_1_51(18) => 
        \DATA_OUT_1_51[18]\, DATA_IN_1_51(17) => 
        \DATA_OUT_1_51[17]\, DATA_IN_1_51(16) => 
        \DATA_OUT_1_51[16]\, DATA_IN_1_51(15) => 
        \DATA_OUT_1_51[15]\, DATA_IN_1_51(14) => 
        \DATA_OUT_1_51[14]\, DATA_IN_1_51(13) => 
        \DATA_OUT_1_51[13]\, DATA_IN_1_51(12) => 
        \DATA_OUT_1_51[12]\, DATA_IN_1_51(11) => 
        \DATA_OUT_1_51[11]\, DATA_IN_1_51(10) => 
        \DATA_OUT_1_51[10]\, DATA_IN_1_51(9) => 
        \DATA_OUT_1_51[9]\, DATA_IN_1_51(8) => \DATA_OUT_1_51[8]\, 
        DATA_IN_1_51(7) => \DATA_OUT_1_51[7]\, DATA_IN_1_51(6)
         => \DATA_OUT_1_51[6]\, DATA_IN_1_51(5) => 
        \DATA_OUT_1_51[5]\, DATA_IN_1_51(4) => \DATA_OUT_1_51[4]\, 
        DATA_IN_1_51(3) => \DATA_OUT_1_51[3]\, DATA_IN_1_51(2)
         => \DATA_OUT_1_51[2]\, DATA_IN_1_51(1) => 
        \DATA_OUT_1_51[1]\, DATA_IN_1_51(0) => \DATA_OUT_1_51[0]\, 
        DATA_OUT_0_0(25) => \DATA_OR_0_3[25]\, DATA_OUT_0_0(24)
         => \DATA_OR_0_3[24]\, DATA_OUT_0_0(23) => 
        \DATA_OR_0_3[23]\, DATA_OUT_0_0(22) => \DATA_OR_0_3[22]\, 
        DATA_OUT_0_0(21) => \DATA_OR_0_3[21]\, DATA_OUT_0_0(20)
         => \DATA_OR_0_3[20]\, DATA_OUT_0_0(19) => 
        \DATA_OR_0_3[19]\, DATA_OUT_0_0(18) => \DATA_OR_0_3[18]\, 
        DATA_OUT_0_0(17) => \DATA_OR_0_3[17]\, DATA_OUT_0_0(16)
         => \DATA_OR_0_3[16]\, DATA_OUT_0_0(15) => 
        \DATA_OR_0_3[15]\, DATA_OUT_0_0(14) => \DATA_OR_0_3[14]\, 
        DATA_OUT_0_0(13) => \DATA_OR_0_3[13]\, DATA_OUT_0_0(12)
         => \DATA_OR_0_3[12]\, DATA_OUT_0_0(11) => 
        \DATA_OR_0_3[11]\, DATA_OUT_0_0(10) => \DATA_OR_0_3[10]\, 
        DATA_OUT_0_0(9) => \DATA_OR_0_3[9]\, DATA_OUT_0_0(8) => 
        \DATA_OR_0_3[8]\, DATA_OUT_0_0(7) => \DATA_OR_0_3[7]\, 
        DATA_OUT_0_0(6) => \DATA_OR_0_3[6]\, DATA_OUT_0_0(5) => 
        \DATA_OR_0_3[5]\, DATA_OUT_0_0(4) => \DATA_OR_0_3[4]\, 
        DATA_OUT_0_0(3) => \DATA_OR_0_3[3]\, DATA_OUT_0_0(2) => 
        \DATA_OR_0_3[2]\, DATA_OUT_0_0(1) => \DATA_OR_0_3[1]\, 
        DATA_OUT_0_0(0) => \DATA_OR_0_3[0]\, DATA_OUT_0_1(25) => 
        \DATA_OR_0_0[25]\, DATA_OUT_0_1(24) => \DATA_OR_0_0[24]\, 
        DATA_OUT_0_1(23) => \DATA_OR_0_0[23]\, DATA_OUT_0_1(22)
         => \DATA_OR_0_0[22]\, DATA_OUT_0_1(21) => 
        \DATA_OR_0_0[21]\, DATA_OUT_0_1(20) => \DATA_OR_0_0[20]\, 
        DATA_OUT_0_1(19) => \DATA_OR_0_0[19]\, DATA_OUT_0_1(18)
         => \DATA_OR_0_0[18]\, DATA_OUT_0_1(17) => 
        \DATA_OR_0_0[17]\, DATA_OUT_0_1(16) => \DATA_OR_0_0[16]\, 
        DATA_OUT_0_1(15) => \DATA_OR_0_0[15]\, DATA_OUT_0_1(14)
         => \DATA_OR_0_0[14]\, DATA_OUT_0_1(13) => 
        \DATA_OR_0_0[13]\, DATA_OUT_0_1(12) => \DATA_OR_0_0[12]\, 
        DATA_OUT_0_1(11) => \DATA_OR_0_0[11]\, DATA_OUT_0_1(10)
         => \DATA_OR_0_0[10]\, DATA_OUT_0_1(9) => 
        \DATA_OR_0_0[9]\, DATA_OUT_0_1(8) => \DATA_OR_0_0[8]\, 
        DATA_OUT_0_1(7) => \DATA_OR_0_0[7]\, DATA_OUT_0_1(6) => 
        \DATA_OR_0_0[6]\, DATA_OUT_0_1(5) => \DATA_OR_0_0[5]\, 
        DATA_OUT_0_1(4) => \DATA_OR_0_0[4]\, DATA_OUT_0_1(3) => 
        \DATA_OR_0_0[3]\, DATA_OUT_0_1(2) => \DATA_OR_0_0[2]\, 
        DATA_OUT_0_1(1) => \DATA_OR_0_0[1]\, DATA_OUT_0_1(0) => 
        \DATA_OR_0_0[0]\, DATA_OUT_0_2(25) => \DATA_OR_0_1[25]\, 
        DATA_OUT_0_2(24) => \DATA_OR_0_1[24]\, DATA_OUT_0_2(23)
         => \DATA_OR_0_1[23]\, DATA_OUT_0_2(22) => 
        \DATA_OR_0_1[22]\, DATA_OUT_0_2(21) => \DATA_OR_0_1[21]\, 
        DATA_OUT_0_2(20) => \DATA_OR_0_1[20]\, DATA_OUT_0_2(19)
         => \DATA_OR_0_1[19]\, DATA_OUT_0_2(18) => 
        \DATA_OR_0_1[18]\, DATA_OUT_0_2(17) => \DATA_OR_0_1[17]\, 
        DATA_OUT_0_2(16) => \DATA_OR_0_1[16]\, DATA_OUT_0_2(15)
         => \DATA_OR_0_1[15]\, DATA_OUT_0_2(14) => 
        \DATA_OR_0_1[14]\, DATA_OUT_0_2(13) => \DATA_OR_0_1[13]\, 
        DATA_OUT_0_2(12) => \DATA_OR_0_1[12]\, DATA_OUT_0_2(11)
         => \DATA_OR_0_1[11]\, DATA_OUT_0_2(10) => 
        \DATA_OR_0_1[10]\, DATA_OUT_0_2(9) => \DATA_OR_0_1[9]\, 
        DATA_OUT_0_2(8) => \DATA_OR_0_1[8]\, DATA_OUT_0_2(7) => 
        \DATA_OR_0_1[7]\, DATA_OUT_0_2(6) => \DATA_OR_0_1[6]\, 
        DATA_OUT_0_2(5) => \DATA_OR_0_1[5]\, DATA_OUT_0_2(4) => 
        \DATA_OR_0_1[4]\, DATA_OUT_0_2(3) => \DATA_OR_0_1[3]\, 
        DATA_OUT_0_2(2) => \DATA_OR_0_1[2]\, DATA_OUT_0_2(1) => 
        \DATA_OR_0_1[1]\, DATA_OUT_0_2(0) => \DATA_OR_0_1[0]\, 
        DATA_OUT_0_3(25) => \DATA_OR_0_2[25]\, DATA_OUT_0_3(24)
         => \DATA_OR_0_2[24]\, DATA_OUT_0_3(23) => 
        \DATA_OR_0_2[23]\, DATA_OUT_0_3(22) => \DATA_OR_0_2[22]\, 
        DATA_OUT_0_3(21) => \DATA_OR_0_2[21]\, DATA_OUT_0_3(20)
         => \DATA_OR_0_2[20]\, DATA_OUT_0_3(19) => 
        \DATA_OR_0_2[19]\, DATA_OUT_0_3(18) => \DATA_OR_0_2[18]\, 
        DATA_OUT_0_3(17) => \DATA_OR_0_2[17]\, DATA_OUT_0_3(16)
         => \DATA_OR_0_2[16]\, DATA_OUT_0_3(15) => 
        \DATA_OR_0_2[15]\, DATA_OUT_0_3(14) => \DATA_OR_0_2[14]\, 
        DATA_OUT_0_3(13) => \DATA_OR_0_2[13]\, DATA_OUT_0_3(12)
         => \DATA_OR_0_2[12]\, DATA_OUT_0_3(11) => 
        \DATA_OR_0_2[11]\, DATA_OUT_0_3(10) => \DATA_OR_0_2[10]\, 
        DATA_OUT_0_3(9) => \DATA_OR_0_2[9]\, DATA_OUT_0_3(8) => 
        \DATA_OR_0_2[8]\, DATA_OUT_0_3(7) => \DATA_OR_0_2[7]\, 
        DATA_OUT_0_3(6) => \DATA_OR_0_2[6]\, DATA_OUT_0_3(5) => 
        \DATA_OR_0_2[5]\, DATA_OUT_0_3(4) => \DATA_OR_0_2[4]\, 
        DATA_OUT_0_3(3) => \DATA_OR_0_2[3]\, DATA_OUT_0_3(2) => 
        \DATA_OR_0_2[2]\, DATA_OUT_0_3(1) => \DATA_OR_0_2[1]\, 
        DATA_OUT_0_3(0) => \DATA_OR_0_2[0]\, DATA_OUT_1_0(25) => 
        \DATA_OR_1_0[25]\, DATA_OUT_1_0(24) => \DATA_OR_1_0[24]\, 
        DATA_OUT_1_0(23) => \DATA_OR_1_0[23]\, DATA_OUT_1_0(22)
         => \DATA_OR_1_0[22]\, DATA_OUT_1_0(21) => 
        \DATA_OR_1_0[21]\, DATA_OUT_1_0(20) => \DATA_OR_1_0[20]\, 
        DATA_OUT_1_0(19) => \DATA_OR_1_0[19]\, DATA_OUT_1_0(18)
         => \DATA_OR_1_0[18]\, DATA_OUT_1_0(17) => 
        \DATA_OR_1_0[17]\, DATA_OUT_1_0(16) => \DATA_OR_1_0[16]\, 
        DATA_OUT_1_0(15) => \DATA_OR_1_0[15]\, DATA_OUT_1_0(14)
         => \DATA_OR_1_0[14]\, DATA_OUT_1_0(13) => 
        \DATA_OR_1_0[13]\, DATA_OUT_1_0(12) => \DATA_OR_1_0[12]\, 
        DATA_OUT_1_0(11) => \DATA_OR_1_0[11]\, DATA_OUT_1_0(10)
         => \DATA_OR_1_0[10]\, DATA_OUT_1_0(9) => 
        \DATA_OR_1_0[9]\, DATA_OUT_1_0(8) => \DATA_OR_1_0[8]\, 
        DATA_OUT_1_0(7) => \DATA_OR_1_0[7]\, DATA_OUT_1_0(6) => 
        \DATA_OR_1_0[6]\, DATA_OUT_1_0(5) => \DATA_OR_1_0[5]\, 
        DATA_OUT_1_0(4) => \DATA_OR_1_0[4]\, DATA_OUT_1_0(3) => 
        \DATA_OR_1_0[3]\, DATA_OUT_1_0(2) => \DATA_OR_1_0[2]\, 
        DATA_OUT_1_0(1) => \DATA_OR_1_0[1]\, DATA_OUT_1_0(0) => 
        \DATA_OR_1_0[0]\, DATA_OUT_1_1(25) => \DATA_OR_1_1[25]\, 
        DATA_OUT_1_1(24) => \DATA_OR_1_1[24]\, DATA_OUT_1_1(23)
         => \DATA_OR_1_1[23]\, DATA_OUT_1_1(22) => 
        \DATA_OR_1_1[22]\, DATA_OUT_1_1(21) => \DATA_OR_1_1[21]\, 
        DATA_OUT_1_1(20) => \DATA_OR_1_1[20]\, DATA_OUT_1_1(19)
         => \DATA_OR_1_1[19]\, DATA_OUT_1_1(18) => 
        \DATA_OR_1_1[18]\, DATA_OUT_1_1(17) => \DATA_OR_1_1[17]\, 
        DATA_OUT_1_1(16) => \DATA_OR_1_1[16]\, DATA_OUT_1_1(15)
         => \DATA_OR_1_1[15]\, DATA_OUT_1_1(14) => 
        \DATA_OR_1_1[14]\, DATA_OUT_1_1(13) => \DATA_OR_1_1[13]\, 
        DATA_OUT_1_1(12) => \DATA_OR_1_1[12]\, DATA_OUT_1_1(11)
         => \DATA_OR_1_1[11]\, DATA_OUT_1_1(10) => 
        \DATA_OR_1_1[10]\, DATA_OUT_1_1(9) => \DATA_OR_1_1[9]\, 
        DATA_OUT_1_1(8) => \DATA_OR_1_1[8]\, DATA_OUT_1_1(7) => 
        \DATA_OR_1_1[7]\, DATA_OUT_1_1(6) => \DATA_OR_1_1[6]\, 
        DATA_OUT_1_1(5) => \DATA_OR_1_1[5]\, DATA_OUT_1_1(4) => 
        \DATA_OR_1_1[4]\, DATA_OUT_1_1(3) => \DATA_OR_1_1[3]\, 
        DATA_OUT_1_1(2) => \DATA_OR_1_1[2]\, DATA_OUT_1_1(1) => 
        \DATA_OR_1_1[1]\, DATA_OUT_1_1(0) => \DATA_OR_1_1[0]\, 
        DATA_OUT_1_2(25) => \DATA_OR_1_2[25]\, DATA_OUT_1_2(24)
         => \DATA_OR_1_2[24]\, DATA_OUT_1_2(23) => 
        \DATA_OR_1_2[23]\, DATA_OUT_1_2(22) => \DATA_OR_1_2[22]\, 
        DATA_OUT_1_2(21) => \DATA_OR_1_2[21]\, DATA_OUT_1_2(20)
         => \DATA_OR_1_2[20]\, DATA_OUT_1_2(19) => 
        \DATA_OR_1_2[19]\, DATA_OUT_1_2(18) => \DATA_OR_1_2[18]\, 
        DATA_OUT_1_2(17) => \DATA_OR_1_2[17]\, DATA_OUT_1_2(16)
         => \DATA_OR_1_2[16]\, DATA_OUT_1_2(15) => 
        \DATA_OR_1_2[15]\, DATA_OUT_1_2(14) => \DATA_OR_1_2[14]\, 
        DATA_OUT_1_2(13) => \DATA_OR_1_2[13]\, DATA_OUT_1_2(12)
         => \DATA_OR_1_2[12]\, DATA_OUT_1_2(11) => 
        \DATA_OR_1_2[11]\, DATA_OUT_1_2(10) => \DATA_OR_1_2[10]\, 
        DATA_OUT_1_2(9) => \DATA_OR_1_2[9]\, DATA_OUT_1_2(8) => 
        \DATA_OR_1_2[8]\, DATA_OUT_1_2(7) => \DATA_OR_1_2[7]\, 
        DATA_OUT_1_2(6) => \DATA_OR_1_2[6]\, DATA_OUT_1_2(5) => 
        \DATA_OR_1_2[5]\, DATA_OUT_1_2(4) => \DATA_OR_1_2[4]\, 
        DATA_OUT_1_2(3) => \DATA_OR_1_2[3]\, DATA_OUT_1_2(2) => 
        \DATA_OR_1_2[2]\, DATA_OUT_1_2(1) => \DATA_OR_1_2[1]\, 
        DATA_OUT_1_2(0) => \DATA_OR_1_2[0]\, DATA_OUT_1_3(25) => 
        \DATA_OR_1_3[25]\, DATA_OUT_1_3(24) => \DATA_OR_1_3[24]\, 
        DATA_OUT_1_3(23) => \DATA_OR_1_3[23]\, DATA_OUT_1_3(22)
         => \DATA_OR_1_3[22]\, DATA_OUT_1_3(21) => 
        \DATA_OR_1_3[21]\, DATA_OUT_1_3(20) => \DATA_OR_1_3[20]\, 
        DATA_OUT_1_3(19) => \DATA_OR_1_3[19]\, DATA_OUT_1_3(18)
         => \DATA_OR_1_3[18]\, DATA_OUT_1_3(17) => 
        \DATA_OR_1_3[17]\, DATA_OUT_1_3(16) => \DATA_OR_1_3[16]\, 
        DATA_OUT_1_3(15) => \DATA_OR_1_3[15]\, DATA_OUT_1_3(14)
         => \DATA_OR_1_3[14]\, DATA_OUT_1_3(13) => 
        \DATA_OR_1_3[13]\, DATA_OUT_1_3(12) => \DATA_OR_1_3[12]\, 
        DATA_OUT_1_3(11) => \DATA_OR_1_3[11]\, DATA_OUT_1_3(10)
         => \DATA_OR_1_3[10]\, DATA_OUT_1_3(9) => 
        \DATA_OR_1_3[9]\, DATA_OUT_1_3(8) => \DATA_OR_1_3[8]\, 
        DATA_OUT_1_3(7) => \DATA_OR_1_3[7]\, DATA_OUT_1_3(6) => 
        \DATA_OR_1_3[6]\, DATA_OUT_1_3(5) => \DATA_OR_1_3[5]\, 
        DATA_OUT_1_3(4) => \DATA_OR_1_3[4]\, DATA_OUT_1_3(3) => 
        \DATA_OR_1_3[3]\, DATA_OUT_1_3(2) => \DATA_OR_1_3[2]\, 
        DATA_OUT_1_3(1) => \DATA_OR_1_3[1]\, DATA_OUT_1_3(0) => 
        \DATA_OR_1_3[0]\, DATA_OUT_1_4(25) => \DATA_OR_1_4[25]\, 
        DATA_OUT_1_4(24) => \DATA_OR_1_4[24]\, DATA_OUT_1_4(23)
         => \DATA_OR_1_4[23]\, DATA_OUT_1_4(22) => 
        \DATA_OR_1_4[22]\, DATA_OUT_1_4(21) => \DATA_OR_1_4[21]\, 
        DATA_OUT_1_4(20) => \DATA_OR_1_4[20]\, DATA_OUT_1_4(19)
         => \DATA_OR_1_4[19]\, DATA_OUT_1_4(18) => 
        \DATA_OR_1_4[18]\, DATA_OUT_1_4(17) => \DATA_OR_1_4[17]\, 
        DATA_OUT_1_4(16) => \DATA_OR_1_4[16]\, DATA_OUT_1_4(15)
         => \DATA_OR_1_4[15]\, DATA_OUT_1_4(14) => 
        \DATA_OR_1_4[14]\, DATA_OUT_1_4(13) => \DATA_OR_1_4[13]\, 
        DATA_OUT_1_4(12) => \DATA_OR_1_4[12]\, DATA_OUT_1_4(11)
         => \DATA_OR_1_4[11]\, DATA_OUT_1_4(10) => 
        \DATA_OR_1_4[10]\, DATA_OUT_1_4(9) => \DATA_OR_1_4[9]\, 
        DATA_OUT_1_4(8) => \DATA_OR_1_4[8]\, DATA_OUT_1_4(7) => 
        \DATA_OR_1_4[7]\, DATA_OUT_1_4(6) => \DATA_OR_1_4[6]\, 
        DATA_OUT_1_4(5) => \DATA_OR_1_4[5]\, DATA_OUT_1_4(4) => 
        \DATA_OR_1_4[4]\, DATA_OUT_1_4(3) => \DATA_OR_1_4[3]\, 
        DATA_OUT_1_4(2) => \DATA_OR_1_4[2]\, DATA_OUT_1_4(1) => 
        \DATA_OR_1_4[1]\, DATA_OUT_1_4(0) => \DATA_OR_1_4[0]\, 
        DATA_OUT_1_5(25) => \DATA_OR_1_5[25]\, DATA_OUT_1_5(24)
         => \DATA_OR_1_5[24]\, DATA_OUT_1_5(23) => 
        \DATA_OR_1_5[23]\, DATA_OUT_1_5(22) => \DATA_OR_1_5[22]\, 
        DATA_OUT_1_5(21) => \DATA_OR_1_5[21]\, DATA_OUT_1_5(20)
         => \DATA_OR_1_5[20]\, DATA_OUT_1_5(19) => 
        \DATA_OR_1_5[19]\, DATA_OUT_1_5(18) => \DATA_OR_1_5[18]\, 
        DATA_OUT_1_5(17) => \DATA_OR_1_5[17]\, DATA_OUT_1_5(16)
         => \DATA_OR_1_5[16]\, DATA_OUT_1_5(15) => 
        \DATA_OR_1_5[15]\, DATA_OUT_1_5(14) => \DATA_OR_1_5[14]\, 
        DATA_OUT_1_5(13) => \DATA_OR_1_5[13]\, DATA_OUT_1_5(12)
         => \DATA_OR_1_5[12]\, DATA_OUT_1_5(11) => 
        \DATA_OR_1_5[11]\, DATA_OUT_1_5(10) => \DATA_OR_1_5[10]\, 
        DATA_OUT_1_5(9) => \DATA_OR_1_5[9]\, DATA_OUT_1_5(8) => 
        \DATA_OR_1_5[8]\, DATA_OUT_1_5(7) => \DATA_OR_1_5[7]\, 
        DATA_OUT_1_5(6) => \DATA_OR_1_5[6]\, DATA_OUT_1_5(5) => 
        \DATA_OR_1_5[5]\, DATA_OUT_1_5(4) => \DATA_OR_1_5[4]\, 
        DATA_OUT_1_5(3) => \DATA_OR_1_5[3]\, DATA_OUT_1_5(2) => 
        \DATA_OR_1_5[2]\, DATA_OUT_1_5(1) => \DATA_OR_1_5[1]\, 
        DATA_OUT_1_5(0) => \DATA_OR_1_5[0]\);
    
    Inst_decoder_array : decoder_array
      port map(RST => RST, CLK => CLK, CLR => LATCH, 
        DATA_OUT_0(71) => \WRITE_EN_0[71]\, DATA_OUT_0(70) => 
        \WRITE_EN_0[70]\, DATA_OUT_0(69) => \WRITE_EN_0[69]\, 
        DATA_OUT_0(68) => \WRITE_EN_0[68]\, DATA_OUT_0(67) => 
        \WRITE_EN_0[67]\, DATA_OUT_0(66) => \WRITE_EN_0[66]\, 
        DATA_OUT_0(65) => \WRITE_EN_0[65]\, DATA_OUT_0(64) => 
        \WRITE_EN_0[64]\, DATA_OUT_0(63) => \WRITE_EN_0[63]\, 
        DATA_OUT_0(62) => \WRITE_EN_0[62]\, DATA_OUT_0(61) => 
        \WRITE_EN_0[61]\, DATA_OUT_0(60) => \WRITE_EN_0[60]\, 
        DATA_OUT_0(59) => \WRITE_EN_0[59]\, DATA_OUT_0(58) => 
        \WRITE_EN_0[58]\, DATA_OUT_0(57) => \WRITE_EN_0[57]\, 
        DATA_OUT_0(56) => \WRITE_EN_0[56]\, DATA_OUT_0(55) => 
        \WRITE_EN_0[55]\, DATA_OUT_0(54) => \WRITE_EN_0[54]\, 
        DATA_OUT_0(53) => \WRITE_EN_0[53]\, DATA_OUT_0(52) => 
        \WRITE_EN_0[52]\, DATA_OUT_0(51) => \WRITE_EN_0[51]\, 
        DATA_OUT_0(50) => \WRITE_EN_0[50]\, DATA_OUT_0(49) => 
        \WRITE_EN_0[49]\, DATA_OUT_0(48) => \WRITE_EN_0[48]\, 
        DATA_OUT_0(47) => \WRITE_EN_0[47]\, DATA_OUT_0(46) => 
        \WRITE_EN_0[46]\, DATA_OUT_0(45) => \WRITE_EN_0[45]\, 
        DATA_OUT_0(44) => \WRITE_EN_0[44]\, DATA_OUT_0(43) => 
        \WRITE_EN_0[43]\, DATA_OUT_0(42) => \WRITE_EN_0[42]\, 
        DATA_OUT_0(41) => \WRITE_EN_0[41]\, DATA_OUT_0(40) => 
        \WRITE_EN_0[40]\, DATA_OUT_0(39) => \WRITE_EN_0[39]\, 
        DATA_OUT_0(38) => \WRITE_EN_0[38]\, DATA_OUT_0(37) => 
        \WRITE_EN_0[37]\, DATA_OUT_0(36) => \WRITE_EN_0[36]\, 
        DATA_OUT_0(35) => \WRITE_EN_0[35]\, DATA_OUT_0(34) => 
        \WRITE_EN_0[34]\, DATA_OUT_0(33) => \WRITE_EN_0[33]\, 
        DATA_OUT_0(32) => \WRITE_EN_0[32]\, DATA_OUT_0(31) => 
        \WRITE_EN_0[31]\, DATA_OUT_0(30) => \WRITE_EN_0[30]\, 
        DATA_OUT_0(29) => \WRITE_EN_0[29]\, DATA_OUT_0(28) => 
        \WRITE_EN_0[28]\, DATA_OUT_0(27) => \WRITE_EN_0[27]\, 
        DATA_OUT_0(26) => \WRITE_EN_0[26]\, DATA_OUT_0(25) => 
        \WRITE_EN_0[25]\, DATA_OUT_0(24) => \WRITE_EN_0[24]\, 
        DATA_OUT_0(23) => \WRITE_EN_0[23]\, DATA_OUT_0(22) => 
        \WRITE_EN_0[22]\, DATA_OUT_0(21) => \WRITE_EN_0[21]\, 
        DATA_OUT_0(20) => \WRITE_EN_0[20]\, DATA_OUT_0(19) => 
        \WRITE_EN_0[19]\, DATA_OUT_0(18) => \WRITE_EN_0[18]\, 
        DATA_OUT_0(17) => \WRITE_EN_0[17]\, DATA_OUT_0(16) => 
        \WRITE_EN_0[16]\, DATA_OUT_0(15) => \WRITE_EN_0[15]\, 
        DATA_OUT_0(14) => \WRITE_EN_0[14]\, DATA_OUT_0(13) => 
        \WRITE_EN_0[13]\, DATA_OUT_0(12) => \WRITE_EN_0[12]\, 
        DATA_OUT_0(11) => \WRITE_EN_0[11]\, DATA_OUT_0(10) => 
        \WRITE_EN_0[10]\, DATA_OUT_0(9) => \WRITE_EN_0[9]\, 
        DATA_OUT_0(8) => \WRITE_EN_0[8]\, DATA_OUT_0(7) => 
        \WRITE_EN_0[7]\, DATA_OUT_0(6) => \WRITE_EN_0[6]\, 
        DATA_OUT_0(5) => \WRITE_EN_0[5]\, DATA_OUT_0(4) => 
        \WRITE_EN_0[4]\, DATA_OUT_0(3) => \WRITE_EN_0[3]\, 
        DATA_OUT_0(2) => \WRITE_EN_0[2]\, DATA_OUT_0(1) => 
        \WRITE_EN_0[1]\, DATA_OUT_0(0) => \WRITE_EN_0[0]\, 
        DATA_OUT_1(103) => \WRITE_EN_1[103]\, DATA_OUT_1(102) => 
        \WRITE_EN_1[102]\, DATA_OUT_1(101) => \WRITE_EN_1[101]\, 
        DATA_OUT_1(100) => \WRITE_EN_1[100]\, DATA_OUT_1(99) => 
        \WRITE_EN_1[99]\, DATA_OUT_1(98) => \WRITE_EN_1[98]\, 
        DATA_OUT_1(97) => \WRITE_EN_1[97]\, DATA_OUT_1(96) => 
        \WRITE_EN_1[96]\, DATA_OUT_1(95) => \WRITE_EN_1[95]\, 
        DATA_OUT_1(94) => \WRITE_EN_1[94]\, DATA_OUT_1(93) => 
        \WRITE_EN_1[93]\, DATA_OUT_1(92) => \WRITE_EN_1[92]\, 
        DATA_OUT_1(91) => \WRITE_EN_1[91]\, DATA_OUT_1(90) => 
        \WRITE_EN_1[90]\, DATA_OUT_1(89) => \WRITE_EN_1[89]\, 
        DATA_OUT_1(88) => \WRITE_EN_1[88]\, DATA_OUT_1(87) => 
        \WRITE_EN_1[87]\, DATA_OUT_1(86) => \WRITE_EN_1[86]\, 
        DATA_OUT_1(85) => \WRITE_EN_1[85]\, DATA_OUT_1(84) => 
        \WRITE_EN_1[84]\, DATA_OUT_1(83) => \WRITE_EN_1[83]\, 
        DATA_OUT_1(82) => \WRITE_EN_1[82]\, DATA_OUT_1(81) => 
        \WRITE_EN_1[81]\, DATA_OUT_1(80) => \WRITE_EN_1[80]\, 
        DATA_OUT_1(79) => \WRITE_EN_1[79]\, DATA_OUT_1(78) => 
        \WRITE_EN_1[78]\, DATA_OUT_1(77) => \WRITE_EN_1[77]\, 
        DATA_OUT_1(76) => \WRITE_EN_1[76]\, DATA_OUT_1(75) => 
        \WRITE_EN_1[75]\, DATA_OUT_1(74) => \WRITE_EN_1[74]\, 
        DATA_OUT_1(73) => \WRITE_EN_1[73]\, DATA_OUT_1(72) => 
        \WRITE_EN_1[72]\, DATA_OUT_1(71) => \WRITE_EN_1[71]\, 
        DATA_OUT_1(70) => \WRITE_EN_1[70]\, DATA_OUT_1(69) => 
        \WRITE_EN_1[69]\, DATA_OUT_1(68) => \WRITE_EN_1[68]\, 
        DATA_OUT_1(67) => \WRITE_EN_1[67]\, DATA_OUT_1(66) => 
        \WRITE_EN_1[66]\, DATA_OUT_1(65) => \WRITE_EN_1[65]\, 
        DATA_OUT_1(64) => \WRITE_EN_1[64]\, DATA_OUT_1(63) => 
        \WRITE_EN_1[63]\, DATA_OUT_1(62) => \WRITE_EN_1[62]\, 
        DATA_OUT_1(61) => \WRITE_EN_1[61]\, DATA_OUT_1(60) => 
        \WRITE_EN_1[60]\, DATA_OUT_1(59) => \WRITE_EN_1[59]\, 
        DATA_OUT_1(58) => \WRITE_EN_1[58]\, DATA_OUT_1(57) => 
        \WRITE_EN_1[57]\, DATA_OUT_1(56) => \WRITE_EN_1[56]\, 
        DATA_OUT_1(55) => \WRITE_EN_1[55]\, DATA_OUT_1(54) => 
        \WRITE_EN_1[54]\, DATA_OUT_1(53) => \WRITE_EN_1[53]\, 
        DATA_OUT_1(52) => \WRITE_EN_1[52]\, DATA_OUT_1(51) => 
        \WRITE_EN_1[51]\, DATA_OUT_1(50) => \WRITE_EN_1[50]\, 
        DATA_OUT_1(49) => \WRITE_EN_1[49]\, DATA_OUT_1(48) => 
        \WRITE_EN_1[48]\, DATA_OUT_1(47) => \WRITE_EN_1[47]\, 
        DATA_OUT_1(46) => \WRITE_EN_1[46]\, DATA_OUT_1(45) => 
        \WRITE_EN_1[45]\, DATA_OUT_1(44) => \WRITE_EN_1[44]\, 
        DATA_OUT_1(43) => \WRITE_EN_1[43]\, DATA_OUT_1(42) => 
        \WRITE_EN_1[42]\, DATA_OUT_1(41) => \WRITE_EN_1[41]\, 
        DATA_OUT_1(40) => \WRITE_EN_1[40]\, DATA_OUT_1(39) => 
        \WRITE_EN_1[39]\, DATA_OUT_1(38) => \WRITE_EN_1[38]\, 
        DATA_OUT_1(37) => \WRITE_EN_1[37]\, DATA_OUT_1(36) => 
        \WRITE_EN_1[36]\, DATA_OUT_1(35) => \WRITE_EN_1[35]\, 
        DATA_OUT_1(34) => \WRITE_EN_1[34]\, DATA_OUT_1(33) => 
        \WRITE_EN_1[33]\, DATA_OUT_1(32) => \WRITE_EN_1[32]\, 
        DATA_OUT_1(31) => \WRITE_EN_1[31]\, DATA_OUT_1(30) => 
        \WRITE_EN_1[30]\, DATA_OUT_1(29) => \WRITE_EN_1[29]\, 
        DATA_OUT_1(28) => \WRITE_EN_1[28]\, DATA_OUT_1(27) => 
        \WRITE_EN_1[27]\, DATA_OUT_1(26) => \WRITE_EN_1[26]\, 
        DATA_OUT_1(25) => \WRITE_EN_1[25]\, DATA_OUT_1(24) => 
        \WRITE_EN_1[24]\, DATA_OUT_1(23) => \WRITE_EN_1[23]\, 
        DATA_OUT_1(22) => \WRITE_EN_1[22]\, DATA_OUT_1(21) => 
        \WRITE_EN_1[21]\, DATA_OUT_1(20) => \WRITE_EN_1[20]\, 
        DATA_OUT_1(19) => \WRITE_EN_1[19]\, DATA_OUT_1(18) => 
        \WRITE_EN_1[18]\, DATA_OUT_1(17) => \WRITE_EN_1[17]\, 
        DATA_OUT_1(16) => \WRITE_EN_1[16]\, DATA_OUT_1(15) => 
        \WRITE_EN_1[15]\, DATA_OUT_1(14) => \WRITE_EN_1[14]\, 
        DATA_OUT_1(13) => \WRITE_EN_1[13]\, DATA_OUT_1(12) => 
        \WRITE_EN_1[12]\, DATA_OUT_1(11) => \WRITE_EN_1[11]\, 
        DATA_OUT_1(10) => \WRITE_EN_1[10]\, DATA_OUT_1(9) => 
        \WRITE_EN_1[9]\, DATA_OUT_1(8) => \WRITE_EN_1[8]\, 
        DATA_OUT_1(7) => \WRITE_EN_1[7]\, DATA_OUT_1(6) => 
        \WRITE_EN_1[6]\, DATA_OUT_1(5) => \WRITE_EN_1[5]\, 
        DATA_OUT_1(4) => \WRITE_EN_1[4]\, DATA_OUT_1(3) => 
        \WRITE_EN_1[3]\, DATA_OUT_1(2) => \WRITE_EN_1[2]\, 
        DATA_OUT_1(1) => \WRITE_EN_1[1]\, DATA_OUT_1(0) => 
        \WRITE_EN_1[0]\);
    
    Inst_arbiter : output_arbiter
      port map(DATA_IN_0(31) => \GND\, DATA_IN_0(30) => \GND\, 
        DATA_IN_0(29) => \GND\, DATA_IN_0(28) => 
        \DATA_OR_1_0[25]\, DATA_IN_0(27) => \DATA_OR_1_0[18]\, 
        DATA_IN_0(26) => \DATA_OR_1_0[7]\, DATA_IN_0(25) => 
        \DATA_OR_1_0[6]\, DATA_IN_0(24) => \DATA_OR_1_0[5]\, 
        DATA_IN_0(23) => \DATA_OR_1_0[4]\, DATA_IN_0(22) => 
        \DATA_OR_1_0[3]\, DATA_IN_0(21) => \DATA_OR_1_0[2]\, 
        DATA_IN_0(20) => \DATA_OR_1_0[1]\, DATA_IN_0(19) => 
        \DATA_OR_1_0[17]\, DATA_IN_0(18) => \DATA_OR_1_0[16]\, 
        DATA_IN_0(17) => \DATA_OR_1_0[15]\, DATA_IN_0(16) => 
        \DATA_OR_1_0[0]\, DATA_IN_0(15) => \GND\, DATA_IN_0(14)
         => \GND\, DATA_IN_0(13) => \DATA_OR_1_0[24]\, 
        DATA_IN_0(12) => \DATA_OR_1_0[23]\, DATA_IN_0(11) => 
        \DATA_OR_1_0[22]\, DATA_IN_0(10) => \DATA_OR_1_0[21]\, 
        DATA_IN_0(9) => \DATA_OR_1_0[20]\, DATA_IN_0(8) => 
        \DATA_OR_1_0[19]\, DATA_IN_0(7) => \DATA_OR_1_0[14]\, 
        DATA_IN_0(6) => \DATA_OR_1_0[13]\, DATA_IN_0(5) => 
        \DATA_OR_1_0[12]\, DATA_IN_0(4) => \DATA_OR_1_0[11]\, 
        DATA_IN_0(3) => \DATA_OR_1_0[10]\, DATA_IN_0(2) => 
        \DATA_OR_1_0[9]\, DATA_IN_0(1) => \DATA_OR_1_0[8]\, 
        DATA_IN_0(0) => \DATA_OR_1_0[0]\, DATA_IN_1(31) => \GND\, 
        DATA_IN_1(30) => \GND\, DATA_IN_1(29) => \GND\, 
        DATA_IN_1(28) => \DATA_OR_1_1[25]\, DATA_IN_1(27) => 
        \DATA_OR_1_1[18]\, DATA_IN_1(26) => \DATA_OR_1_1[7]\, 
        DATA_IN_1(25) => \DATA_OR_1_1[6]\, DATA_IN_1(24) => 
        \DATA_OR_1_1[5]\, DATA_IN_1(23) => \DATA_OR_1_1[4]\, 
        DATA_IN_1(22) => \DATA_OR_1_1[3]\, DATA_IN_1(21) => 
        \DATA_OR_1_1[2]\, DATA_IN_1(20) => \DATA_OR_1_1[1]\, 
        DATA_IN_1(19) => \DATA_OR_1_1[17]\, DATA_IN_1(18) => 
        \DATA_OR_1_1[16]\, DATA_IN_1(17) => \DATA_OR_1_1[15]\, 
        DATA_IN_1(16) => \DATA_OR_1_1[0]\, DATA_IN_1(15) => \GND\, 
        DATA_IN_1(14) => \GND\, DATA_IN_1(13) => 
        \DATA_OR_1_1[24]\, DATA_IN_1(12) => \DATA_OR_1_1[23]\, 
        DATA_IN_1(11) => \DATA_OR_1_1[22]\, DATA_IN_1(10) => 
        \DATA_OR_1_1[21]\, DATA_IN_1(9) => \DATA_OR_1_1[20]\, 
        DATA_IN_1(8) => \DATA_OR_1_1[19]\, DATA_IN_1(7) => 
        \DATA_OR_1_1[14]\, DATA_IN_1(6) => \DATA_OR_1_1[13]\, 
        DATA_IN_1(5) => \DATA_OR_1_1[12]\, DATA_IN_1(4) => 
        \DATA_OR_1_1[11]\, DATA_IN_1(3) => \DATA_OR_1_1[10]\, 
        DATA_IN_1(2) => \DATA_OR_1_1[9]\, DATA_IN_1(1) => 
        \DATA_OR_1_1[8]\, DATA_IN_1(0) => \DATA_OR_1_1[0]\, 
        DATA_IN_2(31) => \GND\, DATA_IN_2(30) => \GND\, 
        DATA_IN_2(29) => \GND\, DATA_IN_2(28) => 
        \DATA_OR_1_2[25]\, DATA_IN_2(27) => \DATA_OR_1_2[18]\, 
        DATA_IN_2(26) => \DATA_OR_1_2[7]\, DATA_IN_2(25) => 
        \DATA_OR_1_2[6]\, DATA_IN_2(24) => \DATA_OR_1_2[5]\, 
        DATA_IN_2(23) => \DATA_OR_1_2[4]\, DATA_IN_2(22) => 
        \DATA_OR_1_2[3]\, DATA_IN_2(21) => \DATA_OR_1_2[2]\, 
        DATA_IN_2(20) => \DATA_OR_1_2[1]\, DATA_IN_2(19) => 
        \DATA_OR_1_2[17]\, DATA_IN_2(18) => \DATA_OR_1_2[16]\, 
        DATA_IN_2(17) => \DATA_OR_1_2[15]\, DATA_IN_2(16) => 
        \DATA_OR_1_2[0]\, DATA_IN_2(15) => \GND\, DATA_IN_2(14)
         => \GND\, DATA_IN_2(13) => \DATA_OR_1_2[24]\, 
        DATA_IN_2(12) => \DATA_OR_1_2[23]\, DATA_IN_2(11) => 
        \DATA_OR_1_2[22]\, DATA_IN_2(10) => \DATA_OR_1_2[21]\, 
        DATA_IN_2(9) => \DATA_OR_1_2[20]\, DATA_IN_2(8) => 
        \DATA_OR_1_2[19]\, DATA_IN_2(7) => \DATA_OR_1_2[14]\, 
        DATA_IN_2(6) => \DATA_OR_1_2[13]\, DATA_IN_2(5) => 
        \DATA_OR_1_2[12]\, DATA_IN_2(4) => \DATA_OR_1_2[11]\, 
        DATA_IN_2(3) => \DATA_OR_1_2[10]\, DATA_IN_2(2) => 
        \DATA_OR_1_2[9]\, DATA_IN_2(1) => \DATA_OR_1_2[8]\, 
        DATA_IN_2(0) => \DATA_OR_1_2[0]\, DATA_IN_3(31) => \GND\, 
        DATA_IN_3(30) => \GND\, DATA_IN_3(29) => \GND\, 
        DATA_IN_3(28) => \DATA_OR_1_3[25]\, DATA_IN_3(27) => 
        \DATA_OR_1_3[18]\, DATA_IN_3(26) => \DATA_OR_1_3[7]\, 
        DATA_IN_3(25) => \DATA_OR_1_3[6]\, DATA_IN_3(24) => 
        \DATA_OR_1_3[5]\, DATA_IN_3(23) => \DATA_OR_1_3[4]\, 
        DATA_IN_3(22) => \DATA_OR_1_3[3]\, DATA_IN_3(21) => 
        \DATA_OR_1_3[2]\, DATA_IN_3(20) => \DATA_OR_1_3[1]\, 
        DATA_IN_3(19) => \DATA_OR_1_3[17]\, DATA_IN_3(18) => 
        \DATA_OR_1_3[16]\, DATA_IN_3(17) => \DATA_OR_1_3[15]\, 
        DATA_IN_3(16) => \DATA_OR_1_3[0]\, DATA_IN_3(15) => \GND\, 
        DATA_IN_3(14) => \GND\, DATA_IN_3(13) => 
        \DATA_OR_1_3[24]\, DATA_IN_3(12) => \DATA_OR_1_3[23]\, 
        DATA_IN_3(11) => \DATA_OR_1_3[22]\, DATA_IN_3(10) => 
        \DATA_OR_1_3[21]\, DATA_IN_3(9) => \DATA_OR_1_3[20]\, 
        DATA_IN_3(8) => \DATA_OR_1_3[19]\, DATA_IN_3(7) => 
        \DATA_OR_1_3[14]\, DATA_IN_3(6) => \DATA_OR_1_3[13]\, 
        DATA_IN_3(5) => \DATA_OR_1_3[12]\, DATA_IN_3(4) => 
        \DATA_OR_1_3[11]\, DATA_IN_3(3) => \DATA_OR_1_3[10]\, 
        DATA_IN_3(2) => \DATA_OR_1_3[9]\, DATA_IN_3(1) => 
        \DATA_OR_1_3[8]\, DATA_IN_3(0) => \DATA_OR_1_3[0]\, 
        DATA_IN_4(31) => \GND\, DATA_IN_4(30) => \GND\, 
        DATA_IN_4(29) => \GND\, DATA_IN_4(28) => 
        \DATA_OR_1_4[25]\, DATA_IN_4(27) => \DATA_OR_1_4[18]\, 
        DATA_IN_4(26) => \DATA_OR_1_4[7]\, DATA_IN_4(25) => 
        \DATA_OR_1_4[6]\, DATA_IN_4(24) => \DATA_OR_1_4[5]\, 
        DATA_IN_4(23) => \DATA_OR_1_4[4]\, DATA_IN_4(22) => 
        \DATA_OR_1_4[3]\, DATA_IN_4(21) => \DATA_OR_1_4[2]\, 
        DATA_IN_4(20) => \DATA_OR_1_4[1]\, DATA_IN_4(19) => 
        \DATA_OR_1_4[17]\, DATA_IN_4(18) => \DATA_OR_1_4[16]\, 
        DATA_IN_4(17) => \DATA_OR_1_4[15]\, DATA_IN_4(16) => 
        \DATA_OR_1_4[0]\, DATA_IN_4(15) => \GND\, DATA_IN_4(14)
         => \GND\, DATA_IN_4(13) => \DATA_OR_1_4[24]\, 
        DATA_IN_4(12) => \DATA_OR_1_4[23]\, DATA_IN_4(11) => 
        \DATA_OR_1_4[22]\, DATA_IN_4(10) => \DATA_OR_1_4[21]\, 
        DATA_IN_4(9) => \DATA_OR_1_4[20]\, DATA_IN_4(8) => 
        \DATA_OR_1_4[19]\, DATA_IN_4(7) => \DATA_OR_1_4[14]\, 
        DATA_IN_4(6) => \DATA_OR_1_4[13]\, DATA_IN_4(5) => 
        \DATA_OR_1_4[12]\, DATA_IN_4(4) => \DATA_OR_1_4[11]\, 
        DATA_IN_4(3) => \DATA_OR_1_4[10]\, DATA_IN_4(2) => 
        \DATA_OR_1_4[9]\, DATA_IN_4(1) => \DATA_OR_1_4[8]\, 
        DATA_IN_4(0) => \DATA_OR_1_4[0]\, DATA_IN_5(31) => \GND\, 
        DATA_IN_5(30) => \GND\, DATA_IN_5(29) => \GND\, 
        DATA_IN_5(28) => \DATA_OR_1_5[25]\, DATA_IN_5(27) => 
        \DATA_OR_1_5[18]\, DATA_IN_5(26) => \DATA_OR_1_5[7]\, 
        DATA_IN_5(25) => \DATA_OR_1_5[6]\, DATA_IN_5(24) => 
        \DATA_OR_1_5[5]\, DATA_IN_5(23) => \DATA_OR_1_5[4]\, 
        DATA_IN_5(22) => \DATA_OR_1_5[3]\, DATA_IN_5(21) => 
        \DATA_OR_1_5[2]\, DATA_IN_5(20) => \DATA_OR_1_5[1]\, 
        DATA_IN_5(19) => \DATA_OR_1_5[17]\, DATA_IN_5(18) => 
        \DATA_OR_1_5[16]\, DATA_IN_5(17) => \DATA_OR_1_5[15]\, 
        DATA_IN_5(16) => \DATA_OR_1_5[0]\, DATA_IN_5(15) => \GND\, 
        DATA_IN_5(14) => \GND\, DATA_IN_5(13) => 
        \DATA_OR_1_5[24]\, DATA_IN_5(12) => \DATA_OR_1_5[23]\, 
        DATA_IN_5(11) => \DATA_OR_1_5[22]\, DATA_IN_5(10) => 
        \DATA_OR_1_5[21]\, DATA_IN_5(9) => \DATA_OR_1_5[20]\, 
        DATA_IN_5(8) => \DATA_OR_1_5[19]\, DATA_IN_5(7) => 
        \DATA_OR_1_5[14]\, DATA_IN_5(6) => \DATA_OR_1_5[13]\, 
        DATA_IN_5(5) => \DATA_OR_1_5[12]\, DATA_IN_5(4) => 
        \DATA_OR_1_5[11]\, DATA_IN_5(3) => \DATA_OR_1_5[10]\, 
        DATA_IN_5(2) => \DATA_OR_1_5[9]\, DATA_IN_5(1) => 
        \DATA_OR_1_5[8]\, DATA_IN_5(0) => \DATA_OR_1_5[0]\, 
        DATA_IN_6(31) => \GND\, DATA_IN_6(30) => \GND\, 
        DATA_IN_6(29) => \GND\, DATA_IN_6(28) => 
        \DATA_OR_0_0[25]\, DATA_IN_6(27) => \DATA_OR_0_0[18]\, 
        DATA_IN_6(26) => \DATA_OR_0_0[7]\, DATA_IN_6(25) => 
        \DATA_OR_0_0[6]\, DATA_IN_6(24) => \DATA_OR_0_0[5]\, 
        DATA_IN_6(23) => \DATA_OR_0_0[4]\, DATA_IN_6(22) => 
        \DATA_OR_0_0[3]\, DATA_IN_6(21) => \DATA_OR_0_0[2]\, 
        DATA_IN_6(20) => \DATA_OR_0_0[1]\, DATA_IN_6(19) => 
        \DATA_OR_0_0[17]\, DATA_IN_6(18) => \DATA_OR_0_0[16]\, 
        DATA_IN_6(17) => \DATA_OR_0_0[15]\, DATA_IN_6(16) => 
        \DATA_OR_0_0[0]\, DATA_IN_6(15) => \GND\, DATA_IN_6(14)
         => \GND\, DATA_IN_6(13) => \DATA_OR_0_0[24]\, 
        DATA_IN_6(12) => \DATA_OR_0_0[23]\, DATA_IN_6(11) => 
        \DATA_OR_0_0[22]\, DATA_IN_6(10) => \DATA_OR_0_0[21]\, 
        DATA_IN_6(9) => \DATA_OR_0_0[20]\, DATA_IN_6(8) => 
        \DATA_OR_0_0[19]\, DATA_IN_6(7) => \DATA_OR_0_0[14]\, 
        DATA_IN_6(6) => \DATA_OR_0_0[13]\, DATA_IN_6(5) => 
        \DATA_OR_0_0[12]\, DATA_IN_6(4) => \DATA_OR_0_0[11]\, 
        DATA_IN_6(3) => \DATA_OR_0_0[10]\, DATA_IN_6(2) => 
        \DATA_OR_0_0[9]\, DATA_IN_6(1) => \DATA_OR_0_0[8]\, 
        DATA_IN_6(0) => \DATA_OR_0_0[0]\, DATA_IN_7(31) => \GND\, 
        DATA_IN_7(30) => \GND\, DATA_IN_7(29) => \GND\, 
        DATA_IN_7(28) => \DATA_OR_0_1[25]\, DATA_IN_7(27) => 
        \DATA_OR_0_1[18]\, DATA_IN_7(26) => \DATA_OR_0_1[7]\, 
        DATA_IN_7(25) => \DATA_OR_0_1[6]\, DATA_IN_7(24) => 
        \DATA_OR_0_1[5]\, DATA_IN_7(23) => \DATA_OR_0_1[4]\, 
        DATA_IN_7(22) => \DATA_OR_0_1[3]\, DATA_IN_7(21) => 
        \DATA_OR_0_1[2]\, DATA_IN_7(20) => \DATA_OR_0_1[1]\, 
        DATA_IN_7(19) => \DATA_OR_0_1[17]\, DATA_IN_7(18) => 
        \DATA_OR_0_1[16]\, DATA_IN_7(17) => \DATA_OR_0_1[15]\, 
        DATA_IN_7(16) => \DATA_OR_0_1[0]\, DATA_IN_7(15) => \GND\, 
        DATA_IN_7(14) => \GND\, DATA_IN_7(13) => 
        \DATA_OR_0_1[24]\, DATA_IN_7(12) => \DATA_OR_0_1[23]\, 
        DATA_IN_7(11) => \DATA_OR_0_1[22]\, DATA_IN_7(10) => 
        \DATA_OR_0_1[21]\, DATA_IN_7(9) => \DATA_OR_0_1[20]\, 
        DATA_IN_7(8) => \DATA_OR_0_1[19]\, DATA_IN_7(7) => 
        \DATA_OR_0_1[14]\, DATA_IN_7(6) => \DATA_OR_0_1[13]\, 
        DATA_IN_7(5) => \DATA_OR_0_1[12]\, DATA_IN_7(4) => 
        \DATA_OR_0_1[11]\, DATA_IN_7(3) => \DATA_OR_0_1[10]\, 
        DATA_IN_7(2) => \DATA_OR_0_1[9]\, DATA_IN_7(1) => 
        \DATA_OR_0_1[8]\, DATA_IN_7(0) => \DATA_OR_0_1[0]\, 
        DATA_IN_8(31) => \GND\, DATA_IN_8(30) => \GND\, 
        DATA_IN_8(29) => \GND\, DATA_IN_8(28) => 
        \DATA_OR_0_2[25]\, DATA_IN_8(27) => \DATA_OR_0_2[18]\, 
        DATA_IN_8(26) => \DATA_OR_0_2[7]\, DATA_IN_8(25) => 
        \DATA_OR_0_2[6]\, DATA_IN_8(24) => \DATA_OR_0_2[5]\, 
        DATA_IN_8(23) => \DATA_OR_0_2[4]\, DATA_IN_8(22) => 
        \DATA_OR_0_2[3]\, DATA_IN_8(21) => \DATA_OR_0_2[2]\, 
        DATA_IN_8(20) => \DATA_OR_0_2[1]\, DATA_IN_8(19) => 
        \DATA_OR_0_2[17]\, DATA_IN_8(18) => \DATA_OR_0_2[16]\, 
        DATA_IN_8(17) => \DATA_OR_0_2[15]\, DATA_IN_8(16) => 
        \DATA_OR_0_2[0]\, DATA_IN_8(15) => \GND\, DATA_IN_8(14)
         => \GND\, DATA_IN_8(13) => \DATA_OR_0_2[24]\, 
        DATA_IN_8(12) => \DATA_OR_0_2[23]\, DATA_IN_8(11) => 
        \DATA_OR_0_2[22]\, DATA_IN_8(10) => \DATA_OR_0_2[21]\, 
        DATA_IN_8(9) => \DATA_OR_0_2[20]\, DATA_IN_8(8) => 
        \DATA_OR_0_2[19]\, DATA_IN_8(7) => \DATA_OR_0_2[14]\, 
        DATA_IN_8(6) => \DATA_OR_0_2[13]\, DATA_IN_8(5) => 
        \DATA_OR_0_2[12]\, DATA_IN_8(4) => \DATA_OR_0_2[11]\, 
        DATA_IN_8(3) => \DATA_OR_0_2[10]\, DATA_IN_8(2) => 
        \DATA_OR_0_2[9]\, DATA_IN_8(1) => \DATA_OR_0_2[8]\, 
        DATA_IN_8(0) => \DATA_OR_0_2[0]\, DATA_IN_9(31) => \GND\, 
        DATA_IN_9(30) => \GND\, DATA_IN_9(29) => \GND\, 
        DATA_IN_9(28) => \DATA_OR_0_3[25]\, DATA_IN_9(27) => 
        \DATA_OR_0_3[18]\, DATA_IN_9(26) => \DATA_OR_0_3[7]\, 
        DATA_IN_9(25) => \DATA_OR_0_3[6]\, DATA_IN_9(24) => 
        \DATA_OR_0_3[5]\, DATA_IN_9(23) => \DATA_OR_0_3[4]\, 
        DATA_IN_9(22) => \DATA_OR_0_3[3]\, DATA_IN_9(21) => 
        \DATA_OR_0_3[2]\, DATA_IN_9(20) => \DATA_OR_0_3[1]\, 
        DATA_IN_9(19) => \DATA_OR_0_3[17]\, DATA_IN_9(18) => 
        \DATA_OR_0_3[16]\, DATA_IN_9(17) => \DATA_OR_0_3[15]\, 
        DATA_IN_9(16) => \DATA_OR_0_3[0]\, DATA_IN_9(15) => \GND\, 
        DATA_IN_9(14) => \GND\, DATA_IN_9(13) => 
        \DATA_OR_0_3[24]\, DATA_IN_9(12) => \DATA_OR_0_3[23]\, 
        DATA_IN_9(11) => \DATA_OR_0_3[22]\, DATA_IN_9(10) => 
        \DATA_OR_0_3[21]\, DATA_IN_9(9) => \DATA_OR_0_3[20]\, 
        DATA_IN_9(8) => \DATA_OR_0_3[19]\, DATA_IN_9(7) => 
        \DATA_OR_0_3[14]\, DATA_IN_9(6) => \DATA_OR_0_3[13]\, 
        DATA_IN_9(5) => \DATA_OR_0_3[12]\, DATA_IN_9(4) => 
        \DATA_OR_0_3[11]\, DATA_IN_9(3) => \DATA_OR_0_3[10]\, 
        DATA_IN_9(2) => \DATA_OR_0_3[9]\, DATA_IN_9(1) => 
        \DATA_OR_0_3[8]\, DATA_IN_9(0) => \DATA_OR_0_3[0]\, CLK
         => CLK, SEND_DATA_0 => SEND_DATA_0, SEND_DATA_1 => 
        SEND_DATA_1, OUT_CLK => OUT_CLK, DATA_OUT_0(31) => 
        \DATA_OUT_0_tmp[31]\, DATA_OUT_0(30) => 
        \DATA_OUT_0_tmp[30]\, DATA_OUT_0(29) => 
        \DATA_OUT_0_tmp[29]\, DATA_OUT_0(28) => 
        \DATA_OUT_0_tmp[28]\, DATA_OUT_0(27) => 
        \DATA_OUT_0_tmp[27]\, DATA_OUT_0(26) => 
        \DATA_OUT_0_tmp[26]\, DATA_OUT_0(25) => 
        \DATA_OUT_0_tmp[25]\, DATA_OUT_0(24) => 
        \DATA_OUT_0_tmp[24]\, DATA_OUT_0(23) => 
        \DATA_OUT_0_tmp[23]\, DATA_OUT_0(22) => 
        \DATA_OUT_0_tmp[22]\, DATA_OUT_0(21) => 
        \DATA_OUT_0_tmp[21]\, DATA_OUT_0(20) => 
        \DATA_OUT_0_tmp[20]\, DATA_OUT_0(19) => 
        \DATA_OUT_0_tmp[19]\, DATA_OUT_0(18) => 
        \DATA_OUT_0_tmp[18]\, DATA_OUT_0(17) => 
        \DATA_OUT_0_tmp[17]\, DATA_OUT_0(16) => 
        \DATA_OUT_0_tmp[16]\, DATA_OUT_0(15) => 
        \DATA_OUT_0_tmp[15]\, DATA_OUT_0(14) => 
        \DATA_OUT_0_tmp[14]\, DATA_OUT_0(13) => 
        \DATA_OUT_0_tmp[13]\, DATA_OUT_0(12) => 
        \DATA_OUT_0_tmp[12]\, DATA_OUT_0(11) => 
        \DATA_OUT_0_tmp[11]\, DATA_OUT_0(10) => 
        \DATA_OUT_0_tmp[10]\, DATA_OUT_0(9) => 
        \DATA_OUT_0_tmp[9]\, DATA_OUT_0(8) => \DATA_OUT_0_tmp[8]\, 
        DATA_OUT_0(7) => \DATA_OUT_0_tmp[7]\, DATA_OUT_0(6) => 
        \DATA_OUT_0_tmp[6]\, DATA_OUT_0(5) => \DATA_OUT_0_tmp[5]\, 
        DATA_OUT_0(4) => \DATA_OUT_0_tmp[4]\, DATA_OUT_0(3) => 
        \DATA_OUT_0_tmp[3]\, DATA_OUT_0(2) => \DATA_OUT_0_tmp[2]\, 
        DATA_OUT_0(1) => \DATA_OUT_0_tmp[1]\, DATA_OUT_0(0) => 
        \DATA_OUT_0_tmp[0]\, DATA_OUT_1(31) => 
        \DATA_OUT_1_tmp[31]\, DATA_OUT_1(30) => 
        \DATA_OUT_1_tmp[30]\, DATA_OUT_1(29) => 
        \DATA_OUT_1_tmp[29]\, DATA_OUT_1(28) => 
        \DATA_OUT_1_tmp[28]\, DATA_OUT_1(27) => 
        \DATA_OUT_1_tmp[27]\, DATA_OUT_1(26) => 
        \DATA_OUT_1_tmp[26]\, DATA_OUT_1(25) => 
        \DATA_OUT_1_tmp[25]\, DATA_OUT_1(24) => 
        \DATA_OUT_1_tmp[24]\, DATA_OUT_1(23) => 
        \DATA_OUT_1_tmp[23]\, DATA_OUT_1(22) => 
        \DATA_OUT_1_tmp[22]\, DATA_OUT_1(21) => 
        \DATA_OUT_1_tmp[21]\, DATA_OUT_1(20) => 
        \DATA_OUT_1_tmp[20]\, DATA_OUT_1(19) => 
        \DATA_OUT_1_tmp[19]\, DATA_OUT_1(18) => 
        \DATA_OUT_1_tmp[18]\, DATA_OUT_1(17) => 
        \DATA_OUT_1_tmp[17]\, DATA_OUT_1(16) => 
        \DATA_OUT_1_tmp[16]\, DATA_OUT_1(15) => 
        \DATA_OUT_1_tmp[15]\, DATA_OUT_1(14) => 
        \DATA_OUT_1_tmp[14]\, DATA_OUT_1(13) => 
        \DATA_OUT_1_tmp[13]\, DATA_OUT_1(12) => 
        \DATA_OUT_1_tmp[12]\, DATA_OUT_1(11) => 
        \DATA_OUT_1_tmp[11]\, DATA_OUT_1(10) => 
        \DATA_OUT_1_tmp[10]\, DATA_OUT_1(9) => 
        \DATA_OUT_1_tmp[9]\, DATA_OUT_1(8) => \DATA_OUT_1_tmp[8]\, 
        DATA_OUT_1(7) => \DATA_OUT_1_tmp[7]\, DATA_OUT_1(6) => 
        \DATA_OUT_1_tmp[6]\, DATA_OUT_1(5) => \DATA_OUT_1_tmp[5]\, 
        DATA_OUT_1(4) => \DATA_OUT_1_tmp[4]\, DATA_OUT_1(3) => 
        \DATA_OUT_1_tmp[3]\, DATA_OUT_1(2) => \DATA_OUT_1_tmp[2]\, 
        DATA_OUT_1(1) => \DATA_OUT_1_tmp[1]\, DATA_OUT_1(0) => 
        \DATA_OUT_1_tmp[0]\, DATA_OUT_2(31) => 
        \DATA_OUT_2_tmp[31]\, DATA_OUT_2(30) => 
        \DATA_OUT_2_tmp[30]\, DATA_OUT_2(29) => 
        \DATA_OUT_2_tmp[29]\, DATA_OUT_2(28) => 
        \DATA_OUT_2_tmp[28]\, DATA_OUT_2(27) => 
        \DATA_OUT_2_tmp[27]\, DATA_OUT_2(26) => 
        \DATA_OUT_2_tmp[26]\, DATA_OUT_2(25) => 
        \DATA_OUT_2_tmp[25]\, DATA_OUT_2(24) => 
        \DATA_OUT_2_tmp[24]\, DATA_OUT_2(23) => 
        \DATA_OUT_2_tmp[23]\, DATA_OUT_2(22) => 
        \DATA_OUT_2_tmp[22]\, DATA_OUT_2(21) => 
        \DATA_OUT_2_tmp[21]\, DATA_OUT_2(20) => 
        \DATA_OUT_2_tmp[20]\, DATA_OUT_2(19) => 
        \DATA_OUT_2_tmp[19]\, DATA_OUT_2(18) => 
        \DATA_OUT_2_tmp[18]\, DATA_OUT_2(17) => 
        \DATA_OUT_2_tmp[17]\, DATA_OUT_2(16) => 
        \DATA_OUT_2_tmp[16]\, DATA_OUT_2(15) => 
        \DATA_OUT_2_tmp[15]\, DATA_OUT_2(14) => 
        \DATA_OUT_2_tmp[14]\, DATA_OUT_2(13) => 
        \DATA_OUT_2_tmp[13]\, DATA_OUT_2(12) => 
        \DATA_OUT_2_tmp[12]\, DATA_OUT_2(11) => 
        \DATA_OUT_2_tmp[11]\, DATA_OUT_2(10) => 
        \DATA_OUT_2_tmp[10]\, DATA_OUT_2(9) => 
        \DATA_OUT_2_tmp[9]\, DATA_OUT_2(8) => \DATA_OUT_2_tmp[8]\, 
        DATA_OUT_2(7) => \DATA_OUT_2_tmp[7]\, DATA_OUT_2(6) => 
        \DATA_OUT_2_tmp[6]\, DATA_OUT_2(5) => \DATA_OUT_2_tmp[5]\, 
        DATA_OUT_2(4) => \DATA_OUT_2_tmp[4]\, DATA_OUT_2(3) => 
        \DATA_OUT_2_tmp[3]\, DATA_OUT_2(2) => \DATA_OUT_2_tmp[2]\, 
        DATA_OUT_2(1) => \DATA_OUT_2_tmp[1]\, DATA_OUT_2(0) => 
        \DATA_OUT_2_tmp[0]\, DATA_OUT_3(31) => 
        \DATA_OUT_3_tmp[31]\, DATA_OUT_3(30) => 
        \DATA_OUT_3_tmp[30]\, DATA_OUT_3(29) => 
        \DATA_OUT_3_tmp[29]\, DATA_OUT_3(28) => 
        \DATA_OUT_3_tmp[28]\, DATA_OUT_3(27) => 
        \DATA_OUT_3_tmp[27]\, DATA_OUT_3(26) => 
        \DATA_OUT_3_tmp[26]\, DATA_OUT_3(25) => 
        \DATA_OUT_3_tmp[25]\, DATA_OUT_3(24) => 
        \DATA_OUT_3_tmp[24]\, DATA_OUT_3(23) => 
        \DATA_OUT_3_tmp[23]\, DATA_OUT_3(22) => 
        \DATA_OUT_3_tmp[22]\, DATA_OUT_3(21) => 
        \DATA_OUT_3_tmp[21]\, DATA_OUT_3(20) => 
        \DATA_OUT_3_tmp[20]\, DATA_OUT_3(19) => 
        \DATA_OUT_3_tmp[19]\, DATA_OUT_3(18) => 
        \DATA_OUT_3_tmp[18]\, DATA_OUT_3(17) => 
        \DATA_OUT_3_tmp[17]\, DATA_OUT_3(16) => 
        \DATA_OUT_3_tmp[16]\, DATA_OUT_3(15) => 
        \DATA_OUT_3_tmp[15]\, DATA_OUT_3(14) => 
        \DATA_OUT_3_tmp[14]\, DATA_OUT_3(13) => 
        \DATA_OUT_3_tmp[13]\, DATA_OUT_3(12) => 
        \DATA_OUT_3_tmp[12]\, DATA_OUT_3(11) => 
        \DATA_OUT_3_tmp[11]\, DATA_OUT_3(10) => 
        \DATA_OUT_3_tmp[10]\, DATA_OUT_3(9) => 
        \DATA_OUT_3_tmp[9]\, DATA_OUT_3(8) => \DATA_OUT_3_tmp[8]\, 
        DATA_OUT_3(7) => \DATA_OUT_3_tmp[7]\, DATA_OUT_3(6) => 
        \DATA_OUT_3_tmp[6]\, DATA_OUT_3(5) => \DATA_OUT_3_tmp[5]\, 
        DATA_OUT_3(4) => \DATA_OUT_3_tmp[4]\, DATA_OUT_3(3) => 
        \DATA_OUT_3_tmp[3]\, DATA_OUT_3(2) => \DATA_OUT_3_tmp[2]\, 
        DATA_OUT_3(1) => \DATA_OUT_3_tmp[1]\, DATA_OUT_3(0) => 
        \DATA_OUT_3_tmp[0]\, RST => RST);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    Inst_sync_block : sync_block_logic
      port map(RST => RST, CLK => OUT_CLK, DATA_IN_0(31) => 
        \DATA_OUT_0_tmp[31]\, DATA_IN_0(30) => 
        \DATA_OUT_0_tmp[30]\, DATA_IN_0(29) => 
        \DATA_OUT_0_tmp[29]\, DATA_IN_0(28) => 
        \DATA_OUT_0_tmp[28]\, DATA_IN_0(27) => 
        \DATA_OUT_0_tmp[27]\, DATA_IN_0(26) => 
        \DATA_OUT_0_tmp[26]\, DATA_IN_0(25) => 
        \DATA_OUT_0_tmp[25]\, DATA_IN_0(24) => 
        \DATA_OUT_0_tmp[24]\, DATA_IN_0(23) => 
        \DATA_OUT_0_tmp[23]\, DATA_IN_0(22) => 
        \DATA_OUT_0_tmp[22]\, DATA_IN_0(21) => 
        \DATA_OUT_0_tmp[21]\, DATA_IN_0(20) => 
        \DATA_OUT_0_tmp[20]\, DATA_IN_0(19) => 
        \DATA_OUT_0_tmp[19]\, DATA_IN_0(18) => 
        \DATA_OUT_0_tmp[18]\, DATA_IN_0(17) => 
        \DATA_OUT_0_tmp[17]\, DATA_IN_0(16) => 
        \DATA_OUT_0_tmp[16]\, DATA_IN_0(15) => 
        \DATA_OUT_0_tmp[15]\, DATA_IN_0(14) => 
        \DATA_OUT_0_tmp[14]\, DATA_IN_0(13) => 
        \DATA_OUT_0_tmp[13]\, DATA_IN_0(12) => 
        \DATA_OUT_0_tmp[12]\, DATA_IN_0(11) => 
        \DATA_OUT_0_tmp[11]\, DATA_IN_0(10) => 
        \DATA_OUT_0_tmp[10]\, DATA_IN_0(9) => \DATA_OUT_0_tmp[9]\, 
        DATA_IN_0(8) => \DATA_OUT_0_tmp[8]\, DATA_IN_0(7) => 
        \DATA_OUT_0_tmp[7]\, DATA_IN_0(6) => \DATA_OUT_0_tmp[6]\, 
        DATA_IN_0(5) => \DATA_OUT_0_tmp[5]\, DATA_IN_0(4) => 
        \DATA_OUT_0_tmp[4]\, DATA_IN_0(3) => \DATA_OUT_0_tmp[3]\, 
        DATA_IN_0(2) => \DATA_OUT_0_tmp[2]\, DATA_IN_0(1) => 
        \DATA_OUT_0_tmp[1]\, DATA_IN_0(0) => \DATA_OUT_0_tmp[0]\, 
        DATA_IN_1(31) => \DATA_OUT_1_tmp[31]\, DATA_IN_1(30) => 
        \DATA_OUT_1_tmp[30]\, DATA_IN_1(29) => 
        \DATA_OUT_1_tmp[29]\, DATA_IN_1(28) => 
        \DATA_OUT_1_tmp[28]\, DATA_IN_1(27) => 
        \DATA_OUT_1_tmp[27]\, DATA_IN_1(26) => 
        \DATA_OUT_1_tmp[26]\, DATA_IN_1(25) => 
        \DATA_OUT_1_tmp[25]\, DATA_IN_1(24) => 
        \DATA_OUT_1_tmp[24]\, DATA_IN_1(23) => 
        \DATA_OUT_1_tmp[23]\, DATA_IN_1(22) => 
        \DATA_OUT_1_tmp[22]\, DATA_IN_1(21) => 
        \DATA_OUT_1_tmp[21]\, DATA_IN_1(20) => 
        \DATA_OUT_1_tmp[20]\, DATA_IN_1(19) => 
        \DATA_OUT_1_tmp[19]\, DATA_IN_1(18) => 
        \DATA_OUT_1_tmp[18]\, DATA_IN_1(17) => 
        \DATA_OUT_1_tmp[17]\, DATA_IN_1(16) => 
        \DATA_OUT_1_tmp[16]\, DATA_IN_1(15) => 
        \DATA_OUT_1_tmp[15]\, DATA_IN_1(14) => 
        \DATA_OUT_1_tmp[14]\, DATA_IN_1(13) => 
        \DATA_OUT_1_tmp[13]\, DATA_IN_1(12) => 
        \DATA_OUT_1_tmp[12]\, DATA_IN_1(11) => 
        \DATA_OUT_1_tmp[11]\, DATA_IN_1(10) => 
        \DATA_OUT_1_tmp[10]\, DATA_IN_1(9) => \DATA_OUT_1_tmp[9]\, 
        DATA_IN_1(8) => \DATA_OUT_1_tmp[8]\, DATA_IN_1(7) => 
        \DATA_OUT_1_tmp[7]\, DATA_IN_1(6) => \DATA_OUT_1_tmp[6]\, 
        DATA_IN_1(5) => \DATA_OUT_1_tmp[5]\, DATA_IN_1(4) => 
        \DATA_OUT_1_tmp[4]\, DATA_IN_1(3) => \DATA_OUT_1_tmp[3]\, 
        DATA_IN_1(2) => \DATA_OUT_1_tmp[2]\, DATA_IN_1(1) => 
        \DATA_OUT_1_tmp[1]\, DATA_IN_1(0) => \DATA_OUT_1_tmp[0]\, 
        DATA_IN_2(31) => \DATA_OUT_2_tmp[31]\, DATA_IN_2(30) => 
        \DATA_OUT_2_tmp[30]\, DATA_IN_2(29) => 
        \DATA_OUT_2_tmp[29]\, DATA_IN_2(28) => 
        \DATA_OUT_2_tmp[28]\, DATA_IN_2(27) => 
        \DATA_OUT_2_tmp[27]\, DATA_IN_2(26) => 
        \DATA_OUT_2_tmp[26]\, DATA_IN_2(25) => 
        \DATA_OUT_2_tmp[25]\, DATA_IN_2(24) => 
        \DATA_OUT_2_tmp[24]\, DATA_IN_2(23) => 
        \DATA_OUT_2_tmp[23]\, DATA_IN_2(22) => 
        \DATA_OUT_2_tmp[22]\, DATA_IN_2(21) => 
        \DATA_OUT_2_tmp[21]\, DATA_IN_2(20) => 
        \DATA_OUT_2_tmp[20]\, DATA_IN_2(19) => 
        \DATA_OUT_2_tmp[19]\, DATA_IN_2(18) => 
        \DATA_OUT_2_tmp[18]\, DATA_IN_2(17) => 
        \DATA_OUT_2_tmp[17]\, DATA_IN_2(16) => 
        \DATA_OUT_2_tmp[16]\, DATA_IN_2(15) => 
        \DATA_OUT_2_tmp[15]\, DATA_IN_2(14) => 
        \DATA_OUT_2_tmp[14]\, DATA_IN_2(13) => 
        \DATA_OUT_2_tmp[13]\, DATA_IN_2(12) => 
        \DATA_OUT_2_tmp[12]\, DATA_IN_2(11) => 
        \DATA_OUT_2_tmp[11]\, DATA_IN_2(10) => 
        \DATA_OUT_2_tmp[10]\, DATA_IN_2(9) => \DATA_OUT_2_tmp[9]\, 
        DATA_IN_2(8) => \DATA_OUT_2_tmp[8]\, DATA_IN_2(7) => 
        \DATA_OUT_2_tmp[7]\, DATA_IN_2(6) => \DATA_OUT_2_tmp[6]\, 
        DATA_IN_2(5) => \DATA_OUT_2_tmp[5]\, DATA_IN_2(4) => 
        \DATA_OUT_2_tmp[4]\, DATA_IN_2(3) => \DATA_OUT_2_tmp[3]\, 
        DATA_IN_2(2) => \DATA_OUT_2_tmp[2]\, DATA_IN_2(1) => 
        \DATA_OUT_2_tmp[1]\, DATA_IN_2(0) => \DATA_OUT_2_tmp[0]\, 
        DATA_IN_3(31) => \DATA_OUT_3_tmp[31]\, DATA_IN_3(30) => 
        \DATA_OUT_3_tmp[30]\, DATA_IN_3(29) => 
        \DATA_OUT_3_tmp[29]\, DATA_IN_3(28) => 
        \DATA_OUT_3_tmp[28]\, DATA_IN_3(27) => 
        \DATA_OUT_3_tmp[27]\, DATA_IN_3(26) => 
        \DATA_OUT_3_tmp[26]\, DATA_IN_3(25) => 
        \DATA_OUT_3_tmp[25]\, DATA_IN_3(24) => 
        \DATA_OUT_3_tmp[24]\, DATA_IN_3(23) => 
        \DATA_OUT_3_tmp[23]\, DATA_IN_3(22) => 
        \DATA_OUT_3_tmp[22]\, DATA_IN_3(21) => 
        \DATA_OUT_3_tmp[21]\, DATA_IN_3(20) => 
        \DATA_OUT_3_tmp[20]\, DATA_IN_3(19) => 
        \DATA_OUT_3_tmp[19]\, DATA_IN_3(18) => 
        \DATA_OUT_3_tmp[18]\, DATA_IN_3(17) => 
        \DATA_OUT_3_tmp[17]\, DATA_IN_3(16) => 
        \DATA_OUT_3_tmp[16]\, DATA_IN_3(15) => 
        \DATA_OUT_3_tmp[15]\, DATA_IN_3(14) => 
        \DATA_OUT_3_tmp[14]\, DATA_IN_3(13) => 
        \DATA_OUT_3_tmp[13]\, DATA_IN_3(12) => 
        \DATA_OUT_3_tmp[12]\, DATA_IN_3(11) => 
        \DATA_OUT_3_tmp[11]\, DATA_IN_3(10) => 
        \DATA_OUT_3_tmp[10]\, DATA_IN_3(9) => \DATA_OUT_3_tmp[9]\, 
        DATA_IN_3(8) => \DATA_OUT_3_tmp[8]\, DATA_IN_3(7) => 
        \DATA_OUT_3_tmp[7]\, DATA_IN_3(6) => \DATA_OUT_3_tmp[6]\, 
        DATA_IN_3(5) => \DATA_OUT_3_tmp[5]\, DATA_IN_3(4) => 
        \DATA_OUT_3_tmp[4]\, DATA_IN_3(3) => \DATA_OUT_3_tmp[3]\, 
        DATA_IN_3(2) => \DATA_OUT_3_tmp[2]\, DATA_IN_3(1) => 
        \DATA_OUT_3_tmp[1]\, DATA_IN_3(0) => \DATA_OUT_3_tmp[0]\, 
        START => LATCH, LSB(7) => LSB(7), LSB(6) => LSB(6), 
        LSB(5) => LSB(5), LSB(4) => LSB(4), LSB(3) => LSB(3), 
        LSB(2) => LSB(2), LSB(1) => LSB(1), LSB(0) => LSB(0), 
        MSB(7) => MSB(7), MSB(6) => MSB(6), MSB(5) => MSB(5), 
        MSB(4) => MSB(4), MSB(3) => MSB(3), MSB(2) => MSB(2), 
        MSB(1) => MSB(1), MSB(0) => MSB(0), DATA_OUT_0(31) => 
        DATA_OUT_0(31), DATA_OUT_0(30) => DATA_OUT_0(30), 
        DATA_OUT_0(29) => DATA_OUT_0(29), DATA_OUT_0(28) => 
        DATA_OUT_0(28), DATA_OUT_0(27) => DATA_OUT_0(27), 
        DATA_OUT_0(26) => DATA_OUT_0(26), DATA_OUT_0(25) => 
        DATA_OUT_0(25), DATA_OUT_0(24) => DATA_OUT_0(24), 
        DATA_OUT_0(23) => DATA_OUT_0(23), DATA_OUT_0(22) => 
        DATA_OUT_0(22), DATA_OUT_0(21) => DATA_OUT_0(21), 
        DATA_OUT_0(20) => DATA_OUT_0(20), DATA_OUT_0(19) => 
        DATA_OUT_0(19), DATA_OUT_0(18) => DATA_OUT_0(18), 
        DATA_OUT_0(17) => DATA_OUT_0(17), DATA_OUT_0(16) => 
        DATA_OUT_0(16), DATA_OUT_0(15) => DATA_OUT_0(15), 
        DATA_OUT_0(14) => DATA_OUT_0(14), DATA_OUT_0(13) => 
        DATA_OUT_0(13), DATA_OUT_0(12) => DATA_OUT_0(12), 
        DATA_OUT_0(11) => DATA_OUT_0(11), DATA_OUT_0(10) => 
        DATA_OUT_0(10), DATA_OUT_0(9) => DATA_OUT_0(9), 
        DATA_OUT_0(8) => DATA_OUT_0(8), DATA_OUT_0(7) => 
        DATA_OUT_0(7), DATA_OUT_0(6) => DATA_OUT_0(6), 
        DATA_OUT_0(5) => DATA_OUT_0(5), DATA_OUT_0(4) => 
        DATA_OUT_0(4), DATA_OUT_0(3) => DATA_OUT_0(3), 
        DATA_OUT_0(2) => DATA_OUT_0(2), DATA_OUT_0(1) => 
        DATA_OUT_0(1), DATA_OUT_0(0) => DATA_OUT_0(0), 
        DATA_OUT_1(31) => DATA_OUT_1(31), DATA_OUT_1(30) => 
        DATA_OUT_1(30), DATA_OUT_1(29) => DATA_OUT_1(29), 
        DATA_OUT_1(28) => DATA_OUT_1(28), DATA_OUT_1(27) => 
        DATA_OUT_1(27), DATA_OUT_1(26) => DATA_OUT_1(26), 
        DATA_OUT_1(25) => DATA_OUT_1(25), DATA_OUT_1(24) => 
        DATA_OUT_1(24), DATA_OUT_1(23) => DATA_OUT_1(23), 
        DATA_OUT_1(22) => DATA_OUT_1(22), DATA_OUT_1(21) => 
        DATA_OUT_1(21), DATA_OUT_1(20) => DATA_OUT_1(20), 
        DATA_OUT_1(19) => DATA_OUT_1(19), DATA_OUT_1(18) => 
        DATA_OUT_1(18), DATA_OUT_1(17) => DATA_OUT_1(17), 
        DATA_OUT_1(16) => DATA_OUT_1(16), DATA_OUT_1(15) => 
        DATA_OUT_1(15), DATA_OUT_1(14) => DATA_OUT_1(14), 
        DATA_OUT_1(13) => DATA_OUT_1(13), DATA_OUT_1(12) => 
        DATA_OUT_1(12), DATA_OUT_1(11) => DATA_OUT_1(11), 
        DATA_OUT_1(10) => DATA_OUT_1(10), DATA_OUT_1(9) => 
        DATA_OUT_1(9), DATA_OUT_1(8) => DATA_OUT_1(8), 
        DATA_OUT_1(7) => DATA_OUT_1(7), DATA_OUT_1(6) => 
        DATA_OUT_1(6), DATA_OUT_1(5) => DATA_OUT_1(5), 
        DATA_OUT_1(4) => DATA_OUT_1(4), DATA_OUT_1(3) => 
        DATA_OUT_1(3), DATA_OUT_1(2) => DATA_OUT_1(2), 
        DATA_OUT_1(1) => DATA_OUT_1(1), DATA_OUT_1(0) => 
        DATA_OUT_1(0), DATA_OUT_2(31) => DATA_OUT_2(31), 
        DATA_OUT_2(30) => DATA_OUT_2(30), DATA_OUT_2(29) => 
        DATA_OUT_2(29), DATA_OUT_2(28) => DATA_OUT_2(28), 
        DATA_OUT_2(27) => DATA_OUT_2(27), DATA_OUT_2(26) => 
        DATA_OUT_2(26), DATA_OUT_2(25) => DATA_OUT_2(25), 
        DATA_OUT_2(24) => DATA_OUT_2(24), DATA_OUT_2(23) => 
        DATA_OUT_2(23), DATA_OUT_2(22) => DATA_OUT_2(22), 
        DATA_OUT_2(21) => DATA_OUT_2(21), DATA_OUT_2(20) => 
        DATA_OUT_2(20), DATA_OUT_2(19) => DATA_OUT_2(19), 
        DATA_OUT_2(18) => DATA_OUT_2(18), DATA_OUT_2(17) => 
        DATA_OUT_2(17), DATA_OUT_2(16) => DATA_OUT_2(16), 
        DATA_OUT_2(15) => DATA_OUT_2(15), DATA_OUT_2(14) => 
        DATA_OUT_2(14), DATA_OUT_2(13) => DATA_OUT_2(13), 
        DATA_OUT_2(12) => DATA_OUT_2(12), DATA_OUT_2(11) => 
        DATA_OUT_2(11), DATA_OUT_2(10) => DATA_OUT_2(10), 
        DATA_OUT_2(9) => DATA_OUT_2(9), DATA_OUT_2(8) => 
        DATA_OUT_2(8), DATA_OUT_2(7) => DATA_OUT_2(7), 
        DATA_OUT_2(6) => DATA_OUT_2(6), DATA_OUT_2(5) => 
        DATA_OUT_2(5), DATA_OUT_2(4) => DATA_OUT_2(4), 
        DATA_OUT_2(3) => DATA_OUT_2(3), DATA_OUT_2(2) => 
        DATA_OUT_2(2), DATA_OUT_2(1) => DATA_OUT_2(1), 
        DATA_OUT_2(0) => DATA_OUT_2(0), DATA_OUT_3(31) => 
        DATA_OUT_3(31), DATA_OUT_3(30) => DATA_OUT_3(30), 
        DATA_OUT_3(29) => DATA_OUT_3(29), DATA_OUT_3(28) => 
        DATA_OUT_3(28), DATA_OUT_3(27) => DATA_OUT_3(27), 
        DATA_OUT_3(26) => DATA_OUT_3(26), DATA_OUT_3(25) => 
        DATA_OUT_3(25), DATA_OUT_3(24) => DATA_OUT_3(24), 
        DATA_OUT_3(23) => DATA_OUT_3(23), DATA_OUT_3(22) => 
        DATA_OUT_3(22), DATA_OUT_3(21) => DATA_OUT_3(21), 
        DATA_OUT_3(20) => DATA_OUT_3(20), DATA_OUT_3(19) => 
        DATA_OUT_3(19), DATA_OUT_3(18) => DATA_OUT_3(18), 
        DATA_OUT_3(17) => DATA_OUT_3(17), DATA_OUT_3(16) => 
        DATA_OUT_3(16), DATA_OUT_3(15) => DATA_OUT_3(15), 
        DATA_OUT_3(14) => DATA_OUT_3(14), DATA_OUT_3(13) => 
        DATA_OUT_3(13), DATA_OUT_3(12) => DATA_OUT_3(12), 
        DATA_OUT_3(11) => DATA_OUT_3(11), DATA_OUT_3(10) => 
        DATA_OUT_3(10), DATA_OUT_3(9) => DATA_OUT_3(9), 
        DATA_OUT_3(8) => DATA_OUT_3(8), DATA_OUT_3(7) => 
        DATA_OUT_3(7), DATA_OUT_3(6) => DATA_OUT_3(6), 
        DATA_OUT_3(5) => DATA_OUT_3(5), DATA_OUT_3(4) => 
        DATA_OUT_3(4), DATA_OUT_3(3) => DATA_OUT_3(3), 
        DATA_OUT_3(2) => DATA_OUT_3(2), DATA_OUT_3(1) => 
        DATA_OUT_3(1), DATA_OUT_3(0) => DATA_OUT_3(0));
    
    Inst_pf_array : pf_array
      port map(RST => RST, DATA_IN_0(71) => DATA_IN_0(71), 
        DATA_IN_0(70) => DATA_IN_0(70), DATA_IN_0(69) => 
        DATA_IN_0(69), DATA_IN_0(68) => DATA_IN_0(68), 
        DATA_IN_0(67) => DATA_IN_0(67), DATA_IN_0(66) => 
        DATA_IN_0(66), DATA_IN_0(65) => DATA_IN_0(65), 
        DATA_IN_0(64) => DATA_IN_0(64), DATA_IN_0(63) => 
        DATA_IN_0(63), DATA_IN_0(62) => DATA_IN_0(62), 
        DATA_IN_0(61) => DATA_IN_0(61), DATA_IN_0(60) => 
        DATA_IN_0(60), DATA_IN_0(59) => DATA_IN_0(59), 
        DATA_IN_0(58) => DATA_IN_0(58), DATA_IN_0(57) => 
        DATA_IN_0(57), DATA_IN_0(56) => DATA_IN_0(56), 
        DATA_IN_0(55) => DATA_IN_0(55), DATA_IN_0(54) => 
        DATA_IN_0(54), DATA_IN_0(53) => DATA_IN_0(53), 
        DATA_IN_0(52) => DATA_IN_0(52), DATA_IN_0(51) => 
        DATA_IN_0(51), DATA_IN_0(50) => DATA_IN_0(50), 
        DATA_IN_0(49) => DATA_IN_0(49), DATA_IN_0(48) => 
        DATA_IN_0(48), DATA_IN_0(47) => DATA_IN_0(47), 
        DATA_IN_0(46) => DATA_IN_0(46), DATA_IN_0(45) => 
        DATA_IN_0(45), DATA_IN_0(44) => DATA_IN_0(44), 
        DATA_IN_0(43) => DATA_IN_0(43), DATA_IN_0(42) => 
        DATA_IN_0(42), DATA_IN_0(41) => DATA_IN_0(41), 
        DATA_IN_0(40) => DATA_IN_0(40), DATA_IN_0(39) => 
        DATA_IN_0(39), DATA_IN_0(38) => DATA_IN_0(38), 
        DATA_IN_0(37) => DATA_IN_0(37), DATA_IN_0(36) => 
        DATA_IN_0(36), DATA_IN_0(35) => DATA_IN_0(35), 
        DATA_IN_0(34) => DATA_IN_0(34), DATA_IN_0(33) => 
        DATA_IN_0(33), DATA_IN_0(32) => DATA_IN_0(32), 
        DATA_IN_0(31) => DATA_IN_0(31), DATA_IN_0(30) => 
        DATA_IN_0(30), DATA_IN_0(29) => DATA_IN_0(29), 
        DATA_IN_0(28) => DATA_IN_0(28), DATA_IN_0(27) => 
        DATA_IN_0(27), DATA_IN_0(26) => DATA_IN_0(26), 
        DATA_IN_0(25) => DATA_IN_0(25), DATA_IN_0(24) => 
        DATA_IN_0(24), DATA_IN_0(23) => DATA_IN_0(23), 
        DATA_IN_0(22) => DATA_IN_0(22), DATA_IN_0(21) => 
        DATA_IN_0(21), DATA_IN_0(20) => DATA_IN_0(20), 
        DATA_IN_0(19) => DATA_IN_0(19), DATA_IN_0(18) => 
        DATA_IN_0(18), DATA_IN_0(17) => DATA_IN_0(17), 
        DATA_IN_0(16) => DATA_IN_0(16), DATA_IN_0(15) => 
        DATA_IN_0(15), DATA_IN_0(14) => DATA_IN_0(14), 
        DATA_IN_0(13) => DATA_IN_0(13), DATA_IN_0(12) => 
        DATA_IN_0(12), DATA_IN_0(11) => DATA_IN_0(11), 
        DATA_IN_0(10) => DATA_IN_0(10), DATA_IN_0(9) => 
        DATA_IN_0(9), DATA_IN_0(8) => DATA_IN_0(8), DATA_IN_0(7)
         => DATA_IN_0(7), DATA_IN_0(6) => DATA_IN_0(6), 
        DATA_IN_0(5) => DATA_IN_0(5), DATA_IN_0(4) => 
        DATA_IN_0(4), DATA_IN_0(3) => DATA_IN_0(3), DATA_IN_0(2)
         => DATA_IN_0(2), DATA_IN_0(1) => DATA_IN_0(1), 
        DATA_IN_0(0) => DATA_IN_0(0), DATA_IN_1(103) => 
        \DATA_IN_1[103]\, DATA_IN_1(102) => DATA_IN_1(102), 
        DATA_IN_1(101) => DATA_IN_1(101), DATA_IN_1(100) => 
        DATA_IN_1(100), DATA_IN_1(99) => DATA_IN_1(99), 
        DATA_IN_1(98) => DATA_IN_1(98), DATA_IN_1(97) => 
        DATA_IN_1(97), DATA_IN_1(96) => DATA_IN_1(96), 
        DATA_IN_1(95) => DATA_IN_1(95), DATA_IN_1(94) => 
        DATA_IN_1(94), DATA_IN_1(93) => DATA_IN_1(93), 
        DATA_IN_1(92) => DATA_IN_1(92), DATA_IN_1(91) => 
        DATA_IN_1(91), DATA_IN_1(90) => DATA_IN_1(90), 
        DATA_IN_1(89) => DATA_IN_1(89), DATA_IN_1(88) => 
        DATA_IN_1(88), DATA_IN_1(87) => DATA_IN_1(87), 
        DATA_IN_1(86) => DATA_IN_1(86), DATA_IN_1(85) => 
        DATA_IN_1(85), DATA_IN_1(84) => DATA_IN_1(84), 
        DATA_IN_1(83) => DATA_IN_1(83), DATA_IN_1(82) => 
        DATA_IN_1(82), DATA_IN_1(81) => DATA_IN_1(81), 
        DATA_IN_1(80) => DATA_IN_1(80), DATA_IN_1(79) => 
        DATA_IN_1(79), DATA_IN_1(78) => DATA_IN_1(78), 
        DATA_IN_1(77) => DATA_IN_1(77), DATA_IN_1(76) => 
        DATA_IN_1(76), DATA_IN_1(75) => DATA_IN_1(75), 
        DATA_IN_1(74) => DATA_IN_1(74), DATA_IN_1(73) => 
        DATA_IN_1(73), DATA_IN_1(72) => DATA_IN_1(72), 
        DATA_IN_1(71) => DATA_IN_1(71), DATA_IN_1(70) => 
        DATA_IN_1(70), DATA_IN_1(69) => DATA_IN_1(69), 
        DATA_IN_1(68) => DATA_IN_1(68), DATA_IN_1(67) => 
        DATA_IN_1(67), DATA_IN_1(66) => DATA_IN_1(66), 
        DATA_IN_1(65) => DATA_IN_1(65), DATA_IN_1(64) => 
        DATA_IN_1(64), DATA_IN_1(63) => DATA_IN_1(63), 
        DATA_IN_1(62) => DATA_IN_1(62), DATA_IN_1(61) => 
        DATA_IN_1(61), DATA_IN_1(60) => DATA_IN_1(60), 
        DATA_IN_1(59) => DATA_IN_1(59), DATA_IN_1(58) => 
        DATA_IN_1(58), DATA_IN_1(57) => DATA_IN_1(57), 
        DATA_IN_1(56) => DATA_IN_1(56), DATA_IN_1(55) => 
        DATA_IN_1(55), DATA_IN_1(54) => DATA_IN_1(54), 
        DATA_IN_1(53) => DATA_IN_1(53), DATA_IN_1(52) => 
        DATA_IN_1(52), DATA_IN_1(51) => DATA_IN_1(51), 
        DATA_IN_1(50) => DATA_IN_1(50), DATA_IN_1(49) => 
        DATA_IN_1(49), DATA_IN_1(48) => DATA_IN_1(48), 
        DATA_IN_1(47) => DATA_IN_1(47), DATA_IN_1(46) => 
        DATA_IN_1(46), DATA_IN_1(45) => DATA_IN_1(45), 
        DATA_IN_1(44) => DATA_IN_1(44), DATA_IN_1(43) => 
        DATA_IN_1(43), DATA_IN_1(42) => DATA_IN_1(42), 
        DATA_IN_1(41) => DATA_IN_1(41), DATA_IN_1(40) => 
        DATA_IN_1(40), DATA_IN_1(39) => DATA_IN_1(39), 
        DATA_IN_1(38) => DATA_IN_1(38), DATA_IN_1(37) => 
        DATA_IN_1(37), DATA_IN_1(36) => DATA_IN_1(36), 
        DATA_IN_1(35) => DATA_IN_1(35), DATA_IN_1(34) => 
        DATA_IN_1(34), DATA_IN_1(33) => DATA_IN_1(33), 
        DATA_IN_1(32) => DATA_IN_1(32), DATA_IN_1(31) => 
        DATA_IN_1(31), DATA_IN_1(30) => DATA_IN_1(30), 
        DATA_IN_1(29) => DATA_IN_1(29), DATA_IN_1(28) => 
        DATA_IN_1(28), DATA_IN_1(27) => DATA_IN_1(27), 
        DATA_IN_1(26) => DATA_IN_1(26), DATA_IN_1(25) => 
        DATA_IN_1(25), DATA_IN_1(24) => DATA_IN_1(24), 
        DATA_IN_1(23) => DATA_IN_1(23), DATA_IN_1(22) => 
        DATA_IN_1(22), DATA_IN_1(21) => DATA_IN_1(21), 
        DATA_IN_1(20) => DATA_IN_1(20), DATA_IN_1(19) => 
        DATA_IN_1(19), DATA_IN_1(18) => DATA_IN_1(18), 
        DATA_IN_1(17) => DATA_IN_1(17), DATA_IN_1(16) => 
        DATA_IN_1(16), DATA_IN_1(15) => DATA_IN_1(15), 
        DATA_IN_1(14) => DATA_IN_1(14), DATA_IN_1(13) => 
        DATA_IN_1(13), DATA_IN_1(12) => DATA_IN_1(12), 
        DATA_IN_1(11) => DATA_IN_1(11), DATA_IN_1(10) => 
        DATA_IN_1(10), DATA_IN_1(9) => DATA_IN_1(9), DATA_IN_1(8)
         => DATA_IN_1(8), DATA_IN_1(7) => DATA_IN_1(7), 
        DATA_IN_1(6) => DATA_IN_1(6), DATA_IN_1(5) => 
        DATA_IN_1(5), DATA_IN_1(4) => DATA_IN_1(4), DATA_IN_1(3)
         => DATA_IN_1(3), DATA_IN_1(2) => DATA_IN_1(2), 
        DATA_IN_1(1) => DATA_IN_1(1), DATA_IN_1(0) => 
        DATA_IN_1(0), BCO_CLK => BCO_CLK, CLK => CLK, CLK90 => 
        CLK90, LATCH => LATCH, SHIFT_IN => SHIFT_IN, SHIFT_EN => 
        SHIFT_EN, SHIFT_OUT => SHIFT_OUT, DATA_OUT_0(71) => 
        \DATA_OUT_PF_0[71]\, DATA_OUT_0(70) => 
        \DATA_OUT_PF_0[70]\, DATA_OUT_0(69) => 
        \DATA_OUT_PF_0[69]\, DATA_OUT_0(68) => 
        \DATA_OUT_PF_0[68]\, DATA_OUT_0(67) => 
        \DATA_OUT_PF_0[67]\, DATA_OUT_0(66) => 
        \DATA_OUT_PF_0[66]\, DATA_OUT_0(65) => 
        \DATA_OUT_PF_0[65]\, DATA_OUT_0(64) => 
        \DATA_OUT_PF_0[64]\, DATA_OUT_0(63) => 
        \DATA_OUT_PF_0[63]\, DATA_OUT_0(62) => 
        \DATA_OUT_PF_0[62]\, DATA_OUT_0(61) => 
        \DATA_OUT_PF_0[61]\, DATA_OUT_0(60) => 
        \DATA_OUT_PF_0[60]\, DATA_OUT_0(59) => 
        \DATA_OUT_PF_0[59]\, DATA_OUT_0(58) => 
        \DATA_OUT_PF_0[58]\, DATA_OUT_0(57) => 
        \DATA_OUT_PF_0[57]\, DATA_OUT_0(56) => 
        \DATA_OUT_PF_0[56]\, DATA_OUT_0(55) => 
        \DATA_OUT_PF_0[55]\, DATA_OUT_0(54) => 
        \DATA_OUT_PF_0[54]\, DATA_OUT_0(53) => 
        \DATA_OUT_PF_0[53]\, DATA_OUT_0(52) => 
        \DATA_OUT_PF_0[52]\, DATA_OUT_0(51) => 
        \DATA_OUT_PF_0[51]\, DATA_OUT_0(50) => 
        \DATA_OUT_PF_0[50]\, DATA_OUT_0(49) => 
        \DATA_OUT_PF_0[49]\, DATA_OUT_0(48) => 
        \DATA_OUT_PF_0[48]\, DATA_OUT_0(47) => 
        \DATA_OUT_PF_0[47]\, DATA_OUT_0(46) => 
        \DATA_OUT_PF_0[46]\, DATA_OUT_0(45) => 
        \DATA_OUT_PF_0[45]\, DATA_OUT_0(44) => 
        \DATA_OUT_PF_0[44]\, DATA_OUT_0(43) => 
        \DATA_OUT_PF_0[43]\, DATA_OUT_0(42) => 
        \DATA_OUT_PF_0[42]\, DATA_OUT_0(41) => 
        \DATA_OUT_PF_0[41]\, DATA_OUT_0(40) => 
        \DATA_OUT_PF_0[40]\, DATA_OUT_0(39) => 
        \DATA_OUT_PF_0[39]\, DATA_OUT_0(38) => 
        \DATA_OUT_PF_0[38]\, DATA_OUT_0(37) => 
        \DATA_OUT_PF_0[37]\, DATA_OUT_0(36) => 
        \DATA_OUT_PF_0[36]\, DATA_OUT_0(35) => 
        \DATA_OUT_PF_0[35]\, DATA_OUT_0(34) => 
        \DATA_OUT_PF_0[34]\, DATA_OUT_0(33) => 
        \DATA_OUT_PF_0[33]\, DATA_OUT_0(32) => 
        \DATA_OUT_PF_0[32]\, DATA_OUT_0(31) => 
        \DATA_OUT_PF_0[31]\, DATA_OUT_0(30) => 
        \DATA_OUT_PF_0[30]\, DATA_OUT_0(29) => 
        \DATA_OUT_PF_0[29]\, DATA_OUT_0(28) => 
        \DATA_OUT_PF_0[28]\, DATA_OUT_0(27) => 
        \DATA_OUT_PF_0[27]\, DATA_OUT_0(26) => 
        \DATA_OUT_PF_0[26]\, DATA_OUT_0(25) => 
        \DATA_OUT_PF_0[25]\, DATA_OUT_0(24) => 
        \DATA_OUT_PF_0[24]\, DATA_OUT_0(23) => 
        \DATA_OUT_PF_0[23]\, DATA_OUT_0(22) => 
        \DATA_OUT_PF_0[22]\, DATA_OUT_0(21) => 
        \DATA_OUT_PF_0[21]\, DATA_OUT_0(20) => 
        \DATA_OUT_PF_0[20]\, DATA_OUT_0(19) => 
        \DATA_OUT_PF_0[19]\, DATA_OUT_0(18) => 
        \DATA_OUT_PF_0[18]\, DATA_OUT_0(17) => 
        \DATA_OUT_PF_0[17]\, DATA_OUT_0(16) => 
        \DATA_OUT_PF_0[16]\, DATA_OUT_0(15) => 
        \DATA_OUT_PF_0[15]\, DATA_OUT_0(14) => 
        \DATA_OUT_PF_0[14]\, DATA_OUT_0(13) => 
        \DATA_OUT_PF_0[13]\, DATA_OUT_0(12) => 
        \DATA_OUT_PF_0[12]\, DATA_OUT_0(11) => 
        \DATA_OUT_PF_0[11]\, DATA_OUT_0(10) => 
        \DATA_OUT_PF_0[10]\, DATA_OUT_0(9) => \DATA_OUT_PF_0[9]\, 
        DATA_OUT_0(8) => \DATA_OUT_PF_0[8]\, DATA_OUT_0(7) => 
        \DATA_OUT_PF_0[7]\, DATA_OUT_0(6) => \DATA_OUT_PF_0[6]\, 
        DATA_OUT_0(5) => \DATA_OUT_PF_0[5]\, DATA_OUT_0(4) => 
        \DATA_OUT_PF_0[4]\, DATA_OUT_0(3) => \DATA_OUT_PF_0[3]\, 
        DATA_OUT_0(2) => \DATA_OUT_PF_0[2]\, DATA_OUT_0(1) => 
        \DATA_OUT_PF_0[1]\, DATA_OUT_0(0) => \DATA_OUT_PF_0[0]\, 
        DATA_OUT_1(103) => \DATA_OUT_PF_1[103]\, DATA_OUT_1(102)
         => \DATA_OUT_PF_1[102]\, DATA_OUT_1(101) => 
        \DATA_OUT_PF_1[101]\, DATA_OUT_1(100) => 
        \DATA_OUT_PF_1[100]\, DATA_OUT_1(99) => 
        \DATA_OUT_PF_1[99]\, DATA_OUT_1(98) => 
        \DATA_OUT_PF_1[98]\, DATA_OUT_1(97) => 
        \DATA_OUT_PF_1[97]\, DATA_OUT_1(96) => 
        \DATA_OUT_PF_1[96]\, DATA_OUT_1(95) => 
        \DATA_OUT_PF_1[95]\, DATA_OUT_1(94) => 
        \DATA_OUT_PF_1[94]\, DATA_OUT_1(93) => 
        \DATA_OUT_PF_1[93]\, DATA_OUT_1(92) => 
        \DATA_OUT_PF_1[92]\, DATA_OUT_1(91) => 
        \DATA_OUT_PF_1[91]\, DATA_OUT_1(90) => 
        \DATA_OUT_PF_1[90]\, DATA_OUT_1(89) => 
        \DATA_OUT_PF_1[89]\, DATA_OUT_1(88) => 
        \DATA_OUT_PF_1[88]\, DATA_OUT_1(87) => 
        \DATA_OUT_PF_1[87]\, DATA_OUT_1(86) => 
        \DATA_OUT_PF_1[86]\, DATA_OUT_1(85) => 
        \DATA_OUT_PF_1[85]\, DATA_OUT_1(84) => 
        \DATA_OUT_PF_1[84]\, DATA_OUT_1(83) => 
        \DATA_OUT_PF_1[83]\, DATA_OUT_1(82) => 
        \DATA_OUT_PF_1[82]\, DATA_OUT_1(81) => 
        \DATA_OUT_PF_1[81]\, DATA_OUT_1(80) => 
        \DATA_OUT_PF_1[80]\, DATA_OUT_1(79) => 
        \DATA_OUT_PF_1[79]\, DATA_OUT_1(78) => 
        \DATA_OUT_PF_1[78]\, DATA_OUT_1(77) => 
        \DATA_OUT_PF_1[77]\, DATA_OUT_1(76) => 
        \DATA_OUT_PF_1[76]\, DATA_OUT_1(75) => 
        \DATA_OUT_PF_1[75]\, DATA_OUT_1(74) => 
        \DATA_OUT_PF_1[74]\, DATA_OUT_1(73) => 
        \DATA_OUT_PF_1[73]\, DATA_OUT_1(72) => 
        \DATA_OUT_PF_1[72]\, DATA_OUT_1(71) => 
        \DATA_OUT_PF_1[71]\, DATA_OUT_1(70) => 
        \DATA_OUT_PF_1[70]\, DATA_OUT_1(69) => 
        \DATA_OUT_PF_1[69]\, DATA_OUT_1(68) => 
        \DATA_OUT_PF_1[68]\, DATA_OUT_1(67) => 
        \DATA_OUT_PF_1[67]\, DATA_OUT_1(66) => 
        \DATA_OUT_PF_1[66]\, DATA_OUT_1(65) => 
        \DATA_OUT_PF_1[65]\, DATA_OUT_1(64) => 
        \DATA_OUT_PF_1[64]\, DATA_OUT_1(63) => 
        \DATA_OUT_PF_1[63]\, DATA_OUT_1(62) => 
        \DATA_OUT_PF_1[62]\, DATA_OUT_1(61) => 
        \DATA_OUT_PF_1[61]\, DATA_OUT_1(60) => 
        \DATA_OUT_PF_1[60]\, DATA_OUT_1(59) => 
        \DATA_OUT_PF_1[59]\, DATA_OUT_1(58) => 
        \DATA_OUT_PF_1[58]\, DATA_OUT_1(57) => 
        \DATA_OUT_PF_1[57]\, DATA_OUT_1(56) => 
        \DATA_OUT_PF_1[56]\, DATA_OUT_1(55) => 
        \DATA_OUT_PF_1[55]\, DATA_OUT_1(54) => 
        \DATA_OUT_PF_1[54]\, DATA_OUT_1(53) => 
        \DATA_OUT_PF_1[53]\, DATA_OUT_1(52) => 
        \DATA_OUT_PF_1[52]\, DATA_OUT_1(51) => 
        \DATA_OUT_PF_1[51]\, DATA_OUT_1(50) => 
        \DATA_OUT_PF_1[50]\, DATA_OUT_1(49) => 
        \DATA_OUT_PF_1[49]\, DATA_OUT_1(48) => 
        \DATA_OUT_PF_1[48]\, DATA_OUT_1(47) => 
        \DATA_OUT_PF_1[47]\, DATA_OUT_1(46) => 
        \DATA_OUT_PF_1[46]\, DATA_OUT_1(45) => 
        \DATA_OUT_PF_1[45]\, DATA_OUT_1(44) => 
        \DATA_OUT_PF_1[44]\, DATA_OUT_1(43) => 
        \DATA_OUT_PF_1[43]\, DATA_OUT_1(42) => 
        \DATA_OUT_PF_1[42]\, DATA_OUT_1(41) => 
        \DATA_OUT_PF_1[41]\, DATA_OUT_1(40) => 
        \DATA_OUT_PF_1[40]\, DATA_OUT_1(39) => 
        \DATA_OUT_PF_1[39]\, DATA_OUT_1(38) => 
        \DATA_OUT_PF_1[38]\, DATA_OUT_1(37) => 
        \DATA_OUT_PF_1[37]\, DATA_OUT_1(36) => 
        \DATA_OUT_PF_1[36]\, DATA_OUT_1(35) => 
        \DATA_OUT_PF_1[35]\, DATA_OUT_1(34) => 
        \DATA_OUT_PF_1[34]\, DATA_OUT_1(33) => 
        \DATA_OUT_PF_1[33]\, DATA_OUT_1(32) => 
        \DATA_OUT_PF_1[32]\, DATA_OUT_1(31) => 
        \DATA_OUT_PF_1[31]\, DATA_OUT_1(30) => 
        \DATA_OUT_PF_1[30]\, DATA_OUT_1(29) => 
        \DATA_OUT_PF_1[29]\, DATA_OUT_1(28) => 
        \DATA_OUT_PF_1[28]\, DATA_OUT_1(27) => 
        \DATA_OUT_PF_1[27]\, DATA_OUT_1(26) => 
        \DATA_OUT_PF_1[26]\, DATA_OUT_1(25) => 
        \DATA_OUT_PF_1[25]\, DATA_OUT_1(24) => 
        \DATA_OUT_PF_1[24]\, DATA_OUT_1(23) => 
        \DATA_OUT_PF_1[23]\, DATA_OUT_1(22) => 
        \DATA_OUT_PF_1[22]\, DATA_OUT_1(21) => 
        \DATA_OUT_PF_1[21]\, DATA_OUT_1(20) => 
        \DATA_OUT_PF_1[20]\, DATA_OUT_1(19) => 
        \DATA_OUT_PF_1[19]\, DATA_OUT_1(18) => 
        \DATA_OUT_PF_1[18]\, DATA_OUT_1(17) => 
        \DATA_OUT_PF_1[17]\, DATA_OUT_1(16) => 
        \DATA_OUT_PF_1[16]\, DATA_OUT_1(15) => 
        \DATA_OUT_PF_1[15]\, DATA_OUT_1(14) => 
        \DATA_OUT_PF_1[14]\, DATA_OUT_1(13) => 
        \DATA_OUT_PF_1[13]\, DATA_OUT_1(12) => 
        \DATA_OUT_PF_1[12]\, DATA_OUT_1(11) => 
        \DATA_OUT_PF_1[11]\, DATA_OUT_1(10) => 
        \DATA_OUT_PF_1[10]\, DATA_OUT_1(9) => \DATA_OUT_PF_1[9]\, 
        DATA_OUT_1(8) => \DATA_OUT_PF_1[8]\, DATA_OUT_1(7) => 
        \DATA_OUT_PF_1[7]\, DATA_OUT_1(6) => \DATA_OUT_PF_1[6]\, 
        DATA_OUT_1(5) => \DATA_OUT_PF_1[5]\, DATA_OUT_1(4) => 
        \DATA_OUT_PF_1[4]\, DATA_OUT_1(3) => \DATA_OUT_PF_1[3]\, 
        DATA_OUT_1(2) => \DATA_OUT_PF_1[2]\, DATA_OUT_1(1) => 
        \DATA_OUT_PF_1[1]\, DATA_OUT_1(0) => \DATA_OUT_PF_1[0]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    Inst_deser_array : deser_array
      port map(RST => RST, DATA_IN_0(71) => \DATA_OUT_PF_0[71]\, 
        DATA_IN_0(70) => \DATA_OUT_PF_0[70]\, DATA_IN_0(69) => 
        \DATA_OUT_PF_0[69]\, DATA_IN_0(68) => \DATA_OUT_PF_0[68]\, 
        DATA_IN_0(67) => \DATA_OUT_PF_0[67]\, DATA_IN_0(66) => 
        \DATA_OUT_PF_0[66]\, DATA_IN_0(65) => \DATA_OUT_PF_0[65]\, 
        DATA_IN_0(64) => \DATA_OUT_PF_0[64]\, DATA_IN_0(63) => 
        \DATA_OUT_PF_0[63]\, DATA_IN_0(62) => \DATA_OUT_PF_0[62]\, 
        DATA_IN_0(61) => \DATA_OUT_PF_0[61]\, DATA_IN_0(60) => 
        \DATA_OUT_PF_0[60]\, DATA_IN_0(59) => \DATA_OUT_PF_0[59]\, 
        DATA_IN_0(58) => \DATA_OUT_PF_0[58]\, DATA_IN_0(57) => 
        \DATA_OUT_PF_0[57]\, DATA_IN_0(56) => \DATA_OUT_PF_0[56]\, 
        DATA_IN_0(55) => \DATA_OUT_PF_0[55]\, DATA_IN_0(54) => 
        \DATA_OUT_PF_0[54]\, DATA_IN_0(53) => \DATA_OUT_PF_0[53]\, 
        DATA_IN_0(52) => \DATA_OUT_PF_0[52]\, DATA_IN_0(51) => 
        \DATA_OUT_PF_0[51]\, DATA_IN_0(50) => \DATA_OUT_PF_0[50]\, 
        DATA_IN_0(49) => \DATA_OUT_PF_0[49]\, DATA_IN_0(48) => 
        \DATA_OUT_PF_0[48]\, DATA_IN_0(47) => \DATA_OUT_PF_0[47]\, 
        DATA_IN_0(46) => \DATA_OUT_PF_0[46]\, DATA_IN_0(45) => 
        \DATA_OUT_PF_0[45]\, DATA_IN_0(44) => \DATA_OUT_PF_0[44]\, 
        DATA_IN_0(43) => \DATA_OUT_PF_0[43]\, DATA_IN_0(42) => 
        \DATA_OUT_PF_0[42]\, DATA_IN_0(41) => \DATA_OUT_PF_0[41]\, 
        DATA_IN_0(40) => \DATA_OUT_PF_0[40]\, DATA_IN_0(39) => 
        \DATA_OUT_PF_0[39]\, DATA_IN_0(38) => \DATA_OUT_PF_0[38]\, 
        DATA_IN_0(37) => \DATA_OUT_PF_0[37]\, DATA_IN_0(36) => 
        \DATA_OUT_PF_0[36]\, DATA_IN_0(35) => \DATA_OUT_PF_0[35]\, 
        DATA_IN_0(34) => \DATA_OUT_PF_0[34]\, DATA_IN_0(33) => 
        \DATA_OUT_PF_0[33]\, DATA_IN_0(32) => \DATA_OUT_PF_0[32]\, 
        DATA_IN_0(31) => \DATA_OUT_PF_0[31]\, DATA_IN_0(30) => 
        \DATA_OUT_PF_0[30]\, DATA_IN_0(29) => \DATA_OUT_PF_0[29]\, 
        DATA_IN_0(28) => \DATA_OUT_PF_0[28]\, DATA_IN_0(27) => 
        \DATA_OUT_PF_0[27]\, DATA_IN_0(26) => \DATA_OUT_PF_0[26]\, 
        DATA_IN_0(25) => \DATA_OUT_PF_0[25]\, DATA_IN_0(24) => 
        \DATA_OUT_PF_0[24]\, DATA_IN_0(23) => \DATA_OUT_PF_0[23]\, 
        DATA_IN_0(22) => \DATA_OUT_PF_0[22]\, DATA_IN_0(21) => 
        \DATA_OUT_PF_0[21]\, DATA_IN_0(20) => \DATA_OUT_PF_0[20]\, 
        DATA_IN_0(19) => \DATA_OUT_PF_0[19]\, DATA_IN_0(18) => 
        \DATA_OUT_PF_0[18]\, DATA_IN_0(17) => \DATA_OUT_PF_0[17]\, 
        DATA_IN_0(16) => \DATA_OUT_PF_0[16]\, DATA_IN_0(15) => 
        \DATA_OUT_PF_0[15]\, DATA_IN_0(14) => \DATA_OUT_PF_0[14]\, 
        DATA_IN_0(13) => \DATA_OUT_PF_0[13]\, DATA_IN_0(12) => 
        \DATA_OUT_PF_0[12]\, DATA_IN_0(11) => \DATA_OUT_PF_0[11]\, 
        DATA_IN_0(10) => \DATA_OUT_PF_0[10]\, DATA_IN_0(9) => 
        \DATA_OUT_PF_0[9]\, DATA_IN_0(8) => \DATA_OUT_PF_0[8]\, 
        DATA_IN_0(7) => \DATA_OUT_PF_0[7]\, DATA_IN_0(6) => 
        \DATA_OUT_PF_0[6]\, DATA_IN_0(5) => \DATA_OUT_PF_0[5]\, 
        DATA_IN_0(4) => \DATA_OUT_PF_0[4]\, DATA_IN_0(3) => 
        \DATA_OUT_PF_0[3]\, DATA_IN_0(2) => \DATA_OUT_PF_0[2]\, 
        DATA_IN_0(1) => \DATA_OUT_PF_0[1]\, DATA_IN_0(0) => 
        \DATA_OUT_PF_0[0]\, DATA_IN_1(103) => 
        \DATA_OUT_PF_1[103]\, DATA_IN_1(102) => 
        \DATA_OUT_PF_1[102]\, DATA_IN_1(101) => 
        \DATA_OUT_PF_1[101]\, DATA_IN_1(100) => 
        \DATA_OUT_PF_1[100]\, DATA_IN_1(99) => 
        \DATA_OUT_PF_1[99]\, DATA_IN_1(98) => \DATA_OUT_PF_1[98]\, 
        DATA_IN_1(97) => \DATA_OUT_PF_1[97]\, DATA_IN_1(96) => 
        \DATA_OUT_PF_1[96]\, DATA_IN_1(95) => \DATA_OUT_PF_1[95]\, 
        DATA_IN_1(94) => \DATA_OUT_PF_1[94]\, DATA_IN_1(93) => 
        \DATA_OUT_PF_1[93]\, DATA_IN_1(92) => \DATA_OUT_PF_1[92]\, 
        DATA_IN_1(91) => \DATA_OUT_PF_1[91]\, DATA_IN_1(90) => 
        \DATA_OUT_PF_1[90]\, DATA_IN_1(89) => \DATA_OUT_PF_1[89]\, 
        DATA_IN_1(88) => \DATA_OUT_PF_1[88]\, DATA_IN_1(87) => 
        \DATA_OUT_PF_1[87]\, DATA_IN_1(86) => \DATA_OUT_PF_1[86]\, 
        DATA_IN_1(85) => \DATA_OUT_PF_1[85]\, DATA_IN_1(84) => 
        \DATA_OUT_PF_1[84]\, DATA_IN_1(83) => \DATA_OUT_PF_1[83]\, 
        DATA_IN_1(82) => \DATA_OUT_PF_1[82]\, DATA_IN_1(81) => 
        \DATA_OUT_PF_1[81]\, DATA_IN_1(80) => \DATA_OUT_PF_1[80]\, 
        DATA_IN_1(79) => \DATA_OUT_PF_1[79]\, DATA_IN_1(78) => 
        \DATA_OUT_PF_1[78]\, DATA_IN_1(77) => \DATA_OUT_PF_1[77]\, 
        DATA_IN_1(76) => \DATA_OUT_PF_1[76]\, DATA_IN_1(75) => 
        \DATA_OUT_PF_1[75]\, DATA_IN_1(74) => \DATA_OUT_PF_1[74]\, 
        DATA_IN_1(73) => \DATA_OUT_PF_1[73]\, DATA_IN_1(72) => 
        \DATA_OUT_PF_1[72]\, DATA_IN_1(71) => \DATA_OUT_PF_1[71]\, 
        DATA_IN_1(70) => \DATA_OUT_PF_1[70]\, DATA_IN_1(69) => 
        \DATA_OUT_PF_1[69]\, DATA_IN_1(68) => \DATA_OUT_PF_1[68]\, 
        DATA_IN_1(67) => \DATA_OUT_PF_1[67]\, DATA_IN_1(66) => 
        \DATA_OUT_PF_1[66]\, DATA_IN_1(65) => \DATA_OUT_PF_1[65]\, 
        DATA_IN_1(64) => \DATA_OUT_PF_1[64]\, DATA_IN_1(63) => 
        \DATA_OUT_PF_1[63]\, DATA_IN_1(62) => \DATA_OUT_PF_1[62]\, 
        DATA_IN_1(61) => \DATA_OUT_PF_1[61]\, DATA_IN_1(60) => 
        \DATA_OUT_PF_1[60]\, DATA_IN_1(59) => \DATA_OUT_PF_1[59]\, 
        DATA_IN_1(58) => \DATA_OUT_PF_1[58]\, DATA_IN_1(57) => 
        \DATA_OUT_PF_1[57]\, DATA_IN_1(56) => \DATA_OUT_PF_1[56]\, 
        DATA_IN_1(55) => \DATA_OUT_PF_1[55]\, DATA_IN_1(54) => 
        \DATA_OUT_PF_1[54]\, DATA_IN_1(53) => \DATA_OUT_PF_1[53]\, 
        DATA_IN_1(52) => \DATA_OUT_PF_1[52]\, DATA_IN_1(51) => 
        \DATA_OUT_PF_1[51]\, DATA_IN_1(50) => \DATA_OUT_PF_1[50]\, 
        DATA_IN_1(49) => \DATA_OUT_PF_1[49]\, DATA_IN_1(48) => 
        \DATA_OUT_PF_1[48]\, DATA_IN_1(47) => \DATA_OUT_PF_1[47]\, 
        DATA_IN_1(46) => \DATA_OUT_PF_1[46]\, DATA_IN_1(45) => 
        \DATA_OUT_PF_1[45]\, DATA_IN_1(44) => \DATA_OUT_PF_1[44]\, 
        DATA_IN_1(43) => \DATA_OUT_PF_1[43]\, DATA_IN_1(42) => 
        \DATA_OUT_PF_1[42]\, DATA_IN_1(41) => \DATA_OUT_PF_1[41]\, 
        DATA_IN_1(40) => \DATA_OUT_PF_1[40]\, DATA_IN_1(39) => 
        \DATA_OUT_PF_1[39]\, DATA_IN_1(38) => \DATA_OUT_PF_1[38]\, 
        DATA_IN_1(37) => \DATA_OUT_PF_1[37]\, DATA_IN_1(36) => 
        \DATA_OUT_PF_1[36]\, DATA_IN_1(35) => \DATA_OUT_PF_1[35]\, 
        DATA_IN_1(34) => \DATA_OUT_PF_1[34]\, DATA_IN_1(33) => 
        \DATA_OUT_PF_1[33]\, DATA_IN_1(32) => \DATA_OUT_PF_1[32]\, 
        DATA_IN_1(31) => \DATA_OUT_PF_1[31]\, DATA_IN_1(30) => 
        \DATA_OUT_PF_1[30]\, DATA_IN_1(29) => \DATA_OUT_PF_1[29]\, 
        DATA_IN_1(28) => \DATA_OUT_PF_1[28]\, DATA_IN_1(27) => 
        \DATA_OUT_PF_1[27]\, DATA_IN_1(26) => \DATA_OUT_PF_1[26]\, 
        DATA_IN_1(25) => \DATA_OUT_PF_1[25]\, DATA_IN_1(24) => 
        \DATA_OUT_PF_1[24]\, DATA_IN_1(23) => \DATA_OUT_PF_1[23]\, 
        DATA_IN_1(22) => \DATA_OUT_PF_1[22]\, DATA_IN_1(21) => 
        \DATA_OUT_PF_1[21]\, DATA_IN_1(20) => \DATA_OUT_PF_1[20]\, 
        DATA_IN_1(19) => \DATA_OUT_PF_1[19]\, DATA_IN_1(18) => 
        \DATA_OUT_PF_1[18]\, DATA_IN_1(17) => \DATA_OUT_PF_1[17]\, 
        DATA_IN_1(16) => \DATA_OUT_PF_1[16]\, DATA_IN_1(15) => 
        \DATA_OUT_PF_1[15]\, DATA_IN_1(14) => \DATA_OUT_PF_1[14]\, 
        DATA_IN_1(13) => \DATA_OUT_PF_1[13]\, DATA_IN_1(12) => 
        \DATA_OUT_PF_1[12]\, DATA_IN_1(11) => \DATA_OUT_PF_1[11]\, 
        DATA_IN_1(10) => \DATA_OUT_PF_1[10]\, DATA_IN_1(9) => 
        \DATA_OUT_PF_1[9]\, DATA_IN_1(8) => \DATA_OUT_PF_1[8]\, 
        DATA_IN_1(7) => \DATA_OUT_PF_1[7]\, DATA_IN_1(6) => 
        \DATA_OUT_PF_1[6]\, DATA_IN_1(5) => \DATA_OUT_PF_1[5]\, 
        DATA_IN_1(4) => \DATA_OUT_PF_1[4]\, DATA_IN_1(3) => 
        \DATA_OUT_PF_1[3]\, DATA_IN_1(2) => \DATA_OUT_PF_1[2]\, 
        DATA_IN_1(1) => \DATA_OUT_PF_1[1]\, DATA_IN_1(0) => 
        \DATA_OUT_PF_1[0]\, WRITE_EN_0(71) => \WRITE_EN_0[71]\, 
        WRITE_EN_0(70) => \WRITE_EN_0[70]\, WRITE_EN_0(69) => 
        \WRITE_EN_0[69]\, WRITE_EN_0(68) => \WRITE_EN_0[68]\, 
        WRITE_EN_0(67) => \WRITE_EN_0[67]\, WRITE_EN_0(66) => 
        \WRITE_EN_0[66]\, WRITE_EN_0(65) => \WRITE_EN_0[65]\, 
        WRITE_EN_0(64) => \WRITE_EN_0[64]\, WRITE_EN_0(63) => 
        \WRITE_EN_0[63]\, WRITE_EN_0(62) => \WRITE_EN_0[62]\, 
        WRITE_EN_0(61) => \WRITE_EN_0[61]\, WRITE_EN_0(60) => 
        \WRITE_EN_0[60]\, WRITE_EN_0(59) => \WRITE_EN_0[59]\, 
        WRITE_EN_0(58) => \WRITE_EN_0[58]\, WRITE_EN_0(57) => 
        \WRITE_EN_0[57]\, WRITE_EN_0(56) => \WRITE_EN_0[56]\, 
        WRITE_EN_0(55) => \WRITE_EN_0[55]\, WRITE_EN_0(54) => 
        \WRITE_EN_0[54]\, WRITE_EN_0(53) => \WRITE_EN_0[53]\, 
        WRITE_EN_0(52) => \WRITE_EN_0[52]\, WRITE_EN_0(51) => 
        \WRITE_EN_0[51]\, WRITE_EN_0(50) => \WRITE_EN_0[50]\, 
        WRITE_EN_0(49) => \WRITE_EN_0[49]\, WRITE_EN_0(48) => 
        \WRITE_EN_0[48]\, WRITE_EN_0(47) => \WRITE_EN_0[47]\, 
        WRITE_EN_0(46) => \WRITE_EN_0[46]\, WRITE_EN_0(45) => 
        \WRITE_EN_0[45]\, WRITE_EN_0(44) => \WRITE_EN_0[44]\, 
        WRITE_EN_0(43) => \WRITE_EN_0[43]\, WRITE_EN_0(42) => 
        \WRITE_EN_0[42]\, WRITE_EN_0(41) => \WRITE_EN_0[41]\, 
        WRITE_EN_0(40) => \WRITE_EN_0[40]\, WRITE_EN_0(39) => 
        \WRITE_EN_0[39]\, WRITE_EN_0(38) => \WRITE_EN_0[38]\, 
        WRITE_EN_0(37) => \WRITE_EN_0[37]\, WRITE_EN_0(36) => 
        \WRITE_EN_0[36]\, WRITE_EN_0(35) => \WRITE_EN_0[35]\, 
        WRITE_EN_0(34) => \WRITE_EN_0[34]\, WRITE_EN_0(33) => 
        \WRITE_EN_0[33]\, WRITE_EN_0(32) => \WRITE_EN_0[32]\, 
        WRITE_EN_0(31) => \WRITE_EN_0[31]\, WRITE_EN_0(30) => 
        \WRITE_EN_0[30]\, WRITE_EN_0(29) => \WRITE_EN_0[29]\, 
        WRITE_EN_0(28) => \WRITE_EN_0[28]\, WRITE_EN_0(27) => 
        \WRITE_EN_0[27]\, WRITE_EN_0(26) => \WRITE_EN_0[26]\, 
        WRITE_EN_0(25) => \WRITE_EN_0[25]\, WRITE_EN_0(24) => 
        \WRITE_EN_0[24]\, WRITE_EN_0(23) => \WRITE_EN_0[23]\, 
        WRITE_EN_0(22) => \WRITE_EN_0[22]\, WRITE_EN_0(21) => 
        \WRITE_EN_0[21]\, WRITE_EN_0(20) => \WRITE_EN_0[20]\, 
        WRITE_EN_0(19) => \WRITE_EN_0[19]\, WRITE_EN_0(18) => 
        \WRITE_EN_0[18]\, WRITE_EN_0(17) => \WRITE_EN_0[17]\, 
        WRITE_EN_0(16) => \WRITE_EN_0[16]\, WRITE_EN_0(15) => 
        \WRITE_EN_0[15]\, WRITE_EN_0(14) => \WRITE_EN_0[14]\, 
        WRITE_EN_0(13) => \WRITE_EN_0[13]\, WRITE_EN_0(12) => 
        \WRITE_EN_0[12]\, WRITE_EN_0(11) => \WRITE_EN_0[11]\, 
        WRITE_EN_0(10) => \WRITE_EN_0[10]\, WRITE_EN_0(9) => 
        \WRITE_EN_0[9]\, WRITE_EN_0(8) => \WRITE_EN_0[8]\, 
        WRITE_EN_0(7) => \WRITE_EN_0[7]\, WRITE_EN_0(6) => 
        \WRITE_EN_0[6]\, WRITE_EN_0(5) => \WRITE_EN_0[5]\, 
        WRITE_EN_0(4) => \WRITE_EN_0[4]\, WRITE_EN_0(3) => 
        \WRITE_EN_0[3]\, WRITE_EN_0(2) => \WRITE_EN_0[2]\, 
        WRITE_EN_0(1) => \WRITE_EN_0[1]\, WRITE_EN_0(0) => 
        \WRITE_EN_0[0]\, WRITE_EN_1(103) => \WRITE_EN_1[103]\, 
        WRITE_EN_1(102) => \WRITE_EN_1[102]\, WRITE_EN_1(101) => 
        \WRITE_EN_1[101]\, WRITE_EN_1(100) => \WRITE_EN_1[100]\, 
        WRITE_EN_1(99) => \WRITE_EN_1[99]\, WRITE_EN_1(98) => 
        \WRITE_EN_1[98]\, WRITE_EN_1(97) => \WRITE_EN_1[97]\, 
        WRITE_EN_1(96) => \WRITE_EN_1[96]\, WRITE_EN_1(95) => 
        \WRITE_EN_1[95]\, WRITE_EN_1(94) => \WRITE_EN_1[94]\, 
        WRITE_EN_1(93) => \WRITE_EN_1[93]\, WRITE_EN_1(92) => 
        \WRITE_EN_1[92]\, WRITE_EN_1(91) => \WRITE_EN_1[91]\, 
        WRITE_EN_1(90) => \WRITE_EN_1[90]\, WRITE_EN_1(89) => 
        \WRITE_EN_1[89]\, WRITE_EN_1(88) => \WRITE_EN_1[88]\, 
        WRITE_EN_1(87) => \WRITE_EN_1[87]\, WRITE_EN_1(86) => 
        \WRITE_EN_1[86]\, WRITE_EN_1(85) => \WRITE_EN_1[85]\, 
        WRITE_EN_1(84) => \WRITE_EN_1[84]\, WRITE_EN_1(83) => 
        \WRITE_EN_1[83]\, WRITE_EN_1(82) => \WRITE_EN_1[82]\, 
        WRITE_EN_1(81) => \WRITE_EN_1[81]\, WRITE_EN_1(80) => 
        \WRITE_EN_1[80]\, WRITE_EN_1(79) => \WRITE_EN_1[79]\, 
        WRITE_EN_1(78) => \WRITE_EN_1[78]\, WRITE_EN_1(77) => 
        \WRITE_EN_1[77]\, WRITE_EN_1(76) => \WRITE_EN_1[76]\, 
        WRITE_EN_1(75) => \WRITE_EN_1[75]\, WRITE_EN_1(74) => 
        \WRITE_EN_1[74]\, WRITE_EN_1(73) => \WRITE_EN_1[73]\, 
        WRITE_EN_1(72) => \WRITE_EN_1[72]\, WRITE_EN_1(71) => 
        \WRITE_EN_1[71]\, WRITE_EN_1(70) => \WRITE_EN_1[70]\, 
        WRITE_EN_1(69) => \WRITE_EN_1[69]\, WRITE_EN_1(68) => 
        \WRITE_EN_1[68]\, WRITE_EN_1(67) => \WRITE_EN_1[67]\, 
        WRITE_EN_1(66) => \WRITE_EN_1[66]\, WRITE_EN_1(65) => 
        \WRITE_EN_1[65]\, WRITE_EN_1(64) => \WRITE_EN_1[64]\, 
        WRITE_EN_1(63) => \WRITE_EN_1[63]\, WRITE_EN_1(62) => 
        \WRITE_EN_1[62]\, WRITE_EN_1(61) => \WRITE_EN_1[61]\, 
        WRITE_EN_1(60) => \WRITE_EN_1[60]\, WRITE_EN_1(59) => 
        \WRITE_EN_1[59]\, WRITE_EN_1(58) => \WRITE_EN_1[58]\, 
        WRITE_EN_1(57) => \WRITE_EN_1[57]\, WRITE_EN_1(56) => 
        \WRITE_EN_1[56]\, WRITE_EN_1(55) => \WRITE_EN_1[55]\, 
        WRITE_EN_1(54) => \WRITE_EN_1[54]\, WRITE_EN_1(53) => 
        \WRITE_EN_1[53]\, WRITE_EN_1(52) => \WRITE_EN_1[52]\, 
        WRITE_EN_1(51) => \WRITE_EN_1[51]\, WRITE_EN_1(50) => 
        \WRITE_EN_1[50]\, WRITE_EN_1(49) => \WRITE_EN_1[49]\, 
        WRITE_EN_1(48) => \WRITE_EN_1[48]\, WRITE_EN_1(47) => 
        \WRITE_EN_1[47]\, WRITE_EN_1(46) => \WRITE_EN_1[46]\, 
        WRITE_EN_1(45) => \WRITE_EN_1[45]\, WRITE_EN_1(44) => 
        \WRITE_EN_1[44]\, WRITE_EN_1(43) => \WRITE_EN_1[43]\, 
        WRITE_EN_1(42) => \WRITE_EN_1[42]\, WRITE_EN_1(41) => 
        \WRITE_EN_1[41]\, WRITE_EN_1(40) => \WRITE_EN_1[40]\, 
        WRITE_EN_1(39) => \WRITE_EN_1[39]\, WRITE_EN_1(38) => 
        \WRITE_EN_1[38]\, WRITE_EN_1(37) => \WRITE_EN_1[37]\, 
        WRITE_EN_1(36) => \WRITE_EN_1[36]\, WRITE_EN_1(35) => 
        \WRITE_EN_1[35]\, WRITE_EN_1(34) => \WRITE_EN_1[34]\, 
        WRITE_EN_1(33) => \WRITE_EN_1[33]\, WRITE_EN_1(32) => 
        \WRITE_EN_1[32]\, WRITE_EN_1(31) => \WRITE_EN_1[31]\, 
        WRITE_EN_1(30) => \WRITE_EN_1[30]\, WRITE_EN_1(29) => 
        \WRITE_EN_1[29]\, WRITE_EN_1(28) => \WRITE_EN_1[28]\, 
        WRITE_EN_1(27) => \WRITE_EN_1[27]\, WRITE_EN_1(26) => 
        \WRITE_EN_1[26]\, WRITE_EN_1(25) => \WRITE_EN_1[25]\, 
        WRITE_EN_1(24) => \WRITE_EN_1[24]\, WRITE_EN_1(23) => 
        \WRITE_EN_1[23]\, WRITE_EN_1(22) => \WRITE_EN_1[22]\, 
        WRITE_EN_1(21) => \WRITE_EN_1[21]\, WRITE_EN_1(20) => 
        \WRITE_EN_1[20]\, WRITE_EN_1(19) => \WRITE_EN_1[19]\, 
        WRITE_EN_1(18) => \WRITE_EN_1[18]\, WRITE_EN_1(17) => 
        \WRITE_EN_1[17]\, WRITE_EN_1(16) => \WRITE_EN_1[16]\, 
        WRITE_EN_1(15) => \WRITE_EN_1[15]\, WRITE_EN_1(14) => 
        \WRITE_EN_1[14]\, WRITE_EN_1(13) => \WRITE_EN_1[13]\, 
        WRITE_EN_1(12) => \WRITE_EN_1[12]\, WRITE_EN_1(11) => 
        \WRITE_EN_1[11]\, WRITE_EN_1(10) => \WRITE_EN_1[10]\, 
        WRITE_EN_1(9) => \WRITE_EN_1[9]\, WRITE_EN_1(8) => 
        \WRITE_EN_1[8]\, WRITE_EN_1(7) => \WRITE_EN_1[7]\, 
        WRITE_EN_1(6) => \WRITE_EN_1[6]\, WRITE_EN_1(5) => 
        \WRITE_EN_1[5]\, WRITE_EN_1(4) => \WRITE_EN_1[4]\, 
        WRITE_EN_1(3) => \WRITE_EN_1[3]\, WRITE_EN_1(2) => 
        \WRITE_EN_1[2]\, WRITE_EN_1(1) => \WRITE_EN_1[1]\, 
        WRITE_EN_1(0) => \WRITE_EN_1[0]\, CLK => CLK, 
        DATA_OUT_0_0(25) => \DATA_OUT_0_0[25]\, DATA_OUT_0_0(24)
         => \DATA_OUT_0_0[24]\, DATA_OUT_0_0(23) => 
        \DATA_OUT_0_0[23]\, DATA_OUT_0_0(22) => 
        \DATA_OUT_0_0[22]\, DATA_OUT_0_0(21) => 
        \DATA_OUT_0_0[21]\, DATA_OUT_0_0(20) => 
        \DATA_OUT_0_0[20]\, DATA_OUT_0_0(19) => 
        \DATA_OUT_0_0[19]\, DATA_OUT_0_0(18) => 
        \DATA_OUT_0_0[18]\, DATA_OUT_0_0(17) => 
        \DATA_OUT_0_0[17]\, DATA_OUT_0_0(16) => 
        \DATA_OUT_0_0[16]\, DATA_OUT_0_0(15) => 
        \DATA_OUT_0_0[15]\, DATA_OUT_0_0(14) => 
        \DATA_OUT_0_0[14]\, DATA_OUT_0_0(13) => 
        \DATA_OUT_0_0[13]\, DATA_OUT_0_0(12) => 
        \DATA_OUT_0_0[12]\, DATA_OUT_0_0(11) => 
        \DATA_OUT_0_0[11]\, DATA_OUT_0_0(10) => 
        \DATA_OUT_0_0[10]\, DATA_OUT_0_0(9) => \DATA_OUT_0_0[9]\, 
        DATA_OUT_0_0(8) => \DATA_OUT_0_0[8]\, DATA_OUT_0_0(7) => 
        \DATA_OUT_0_0[7]\, DATA_OUT_0_0(6) => \DATA_OUT_0_0[6]\, 
        DATA_OUT_0_0(5) => \DATA_OUT_0_0[5]\, DATA_OUT_0_0(4) => 
        \DATA_OUT_0_0[4]\, DATA_OUT_0_0(3) => \DATA_OUT_0_0[3]\, 
        DATA_OUT_0_0(2) => \DATA_OUT_0_0[2]\, DATA_OUT_0_0(1) => 
        \DATA_OUT_0_0[1]\, DATA_OUT_0_0(0) => \DATA_OUT_0_0[0]\, 
        DATA_OUT_0_1(25) => \DATA_OUT_0_1[25]\, DATA_OUT_0_1(24)
         => \DATA_OUT_0_1[24]\, DATA_OUT_0_1(23) => 
        \DATA_OUT_0_1[23]\, DATA_OUT_0_1(22) => 
        \DATA_OUT_0_1[22]\, DATA_OUT_0_1(21) => 
        \DATA_OUT_0_1[21]\, DATA_OUT_0_1(20) => 
        \DATA_OUT_0_1[20]\, DATA_OUT_0_1(19) => 
        \DATA_OUT_0_1[19]\, DATA_OUT_0_1(18) => 
        \DATA_OUT_0_1[18]\, DATA_OUT_0_1(17) => 
        \DATA_OUT_0_1[17]\, DATA_OUT_0_1(16) => 
        \DATA_OUT_0_1[16]\, DATA_OUT_0_1(15) => 
        \DATA_OUT_0_1[15]\, DATA_OUT_0_1(14) => 
        \DATA_OUT_0_1[14]\, DATA_OUT_0_1(13) => 
        \DATA_OUT_0_1[13]\, DATA_OUT_0_1(12) => 
        \DATA_OUT_0_1[12]\, DATA_OUT_0_1(11) => 
        \DATA_OUT_0_1[11]\, DATA_OUT_0_1(10) => 
        \DATA_OUT_0_1[10]\, DATA_OUT_0_1(9) => \DATA_OUT_0_1[9]\, 
        DATA_OUT_0_1(8) => \DATA_OUT_0_1[8]\, DATA_OUT_0_1(7) => 
        \DATA_OUT_0_1[7]\, DATA_OUT_0_1(6) => \DATA_OUT_0_1[6]\, 
        DATA_OUT_0_1(5) => \DATA_OUT_0_1[5]\, DATA_OUT_0_1(4) => 
        \DATA_OUT_0_1[4]\, DATA_OUT_0_1(3) => \DATA_OUT_0_1[3]\, 
        DATA_OUT_0_1(2) => \DATA_OUT_0_1[2]\, DATA_OUT_0_1(1) => 
        \DATA_OUT_0_1[1]\, DATA_OUT_0_1(0) => \DATA_OUT_0_1[0]\, 
        DATA_OUT_0_2(25) => \DATA_OUT_0_2[25]\, DATA_OUT_0_2(24)
         => \DATA_OUT_0_2[24]\, DATA_OUT_0_2(23) => 
        \DATA_OUT_0_2[23]\, DATA_OUT_0_2(22) => 
        \DATA_OUT_0_2[22]\, DATA_OUT_0_2(21) => 
        \DATA_OUT_0_2[21]\, DATA_OUT_0_2(20) => 
        \DATA_OUT_0_2[20]\, DATA_OUT_0_2(19) => 
        \DATA_OUT_0_2[19]\, DATA_OUT_0_2(18) => 
        \DATA_OUT_0_2[18]\, DATA_OUT_0_2(17) => 
        \DATA_OUT_0_2[17]\, DATA_OUT_0_2(16) => 
        \DATA_OUT_0_2[16]\, DATA_OUT_0_2(15) => 
        \DATA_OUT_0_2[15]\, DATA_OUT_0_2(14) => 
        \DATA_OUT_0_2[14]\, DATA_OUT_0_2(13) => 
        \DATA_OUT_0_2[13]\, DATA_OUT_0_2(12) => 
        \DATA_OUT_0_2[12]\, DATA_OUT_0_2(11) => 
        \DATA_OUT_0_2[11]\, DATA_OUT_0_2(10) => 
        \DATA_OUT_0_2[10]\, DATA_OUT_0_2(9) => \DATA_OUT_0_2[9]\, 
        DATA_OUT_0_2(8) => \DATA_OUT_0_2[8]\, DATA_OUT_0_2(7) => 
        \DATA_OUT_0_2[7]\, DATA_OUT_0_2(6) => \DATA_OUT_0_2[6]\, 
        DATA_OUT_0_2(5) => \DATA_OUT_0_2[5]\, DATA_OUT_0_2(4) => 
        \DATA_OUT_0_2[4]\, DATA_OUT_0_2(3) => \DATA_OUT_0_2[3]\, 
        DATA_OUT_0_2(2) => \DATA_OUT_0_2[2]\, DATA_OUT_0_2(1) => 
        \DATA_OUT_0_2[1]\, DATA_OUT_0_2(0) => \DATA_OUT_0_2[0]\, 
        DATA_OUT_0_3(25) => \DATA_OUT_0_3[25]\, DATA_OUT_0_3(24)
         => \DATA_OUT_0_3[24]\, DATA_OUT_0_3(23) => 
        \DATA_OUT_0_3[23]\, DATA_OUT_0_3(22) => 
        \DATA_OUT_0_3[22]\, DATA_OUT_0_3(21) => 
        \DATA_OUT_0_3[21]\, DATA_OUT_0_3(20) => 
        \DATA_OUT_0_3[20]\, DATA_OUT_0_3(19) => 
        \DATA_OUT_0_3[19]\, DATA_OUT_0_3(18) => 
        \DATA_OUT_0_3[18]\, DATA_OUT_0_3(17) => 
        \DATA_OUT_0_3[17]\, DATA_OUT_0_3(16) => 
        \DATA_OUT_0_3[16]\, DATA_OUT_0_3(15) => 
        \DATA_OUT_0_3[15]\, DATA_OUT_0_3(14) => 
        \DATA_OUT_0_3[14]\, DATA_OUT_0_3(13) => 
        \DATA_OUT_0_3[13]\, DATA_OUT_0_3(12) => 
        \DATA_OUT_0_3[12]\, DATA_OUT_0_3(11) => 
        \DATA_OUT_0_3[11]\, DATA_OUT_0_3(10) => 
        \DATA_OUT_0_3[10]\, DATA_OUT_0_3(9) => \DATA_OUT_0_3[9]\, 
        DATA_OUT_0_3(8) => \DATA_OUT_0_3[8]\, DATA_OUT_0_3(7) => 
        \DATA_OUT_0_3[7]\, DATA_OUT_0_3(6) => \DATA_OUT_0_3[6]\, 
        DATA_OUT_0_3(5) => \DATA_OUT_0_3[5]\, DATA_OUT_0_3(4) => 
        \DATA_OUT_0_3[4]\, DATA_OUT_0_3(3) => \DATA_OUT_0_3[3]\, 
        DATA_OUT_0_3(2) => \DATA_OUT_0_3[2]\, DATA_OUT_0_3(1) => 
        \DATA_OUT_0_3[1]\, DATA_OUT_0_3(0) => \DATA_OUT_0_3[0]\, 
        DATA_OUT_0_4(25) => \DATA_OUT_0_4[25]\, DATA_OUT_0_4(24)
         => \DATA_OUT_0_4[24]\, DATA_OUT_0_4(23) => 
        \DATA_OUT_0_4[23]\, DATA_OUT_0_4(22) => 
        \DATA_OUT_0_4[22]\, DATA_OUT_0_4(21) => 
        \DATA_OUT_0_4[21]\, DATA_OUT_0_4(20) => 
        \DATA_OUT_0_4[20]\, DATA_OUT_0_4(19) => 
        \DATA_OUT_0_4[19]\, DATA_OUT_0_4(18) => 
        \DATA_OUT_0_4[18]\, DATA_OUT_0_4(17) => 
        \DATA_OUT_0_4[17]\, DATA_OUT_0_4(16) => 
        \DATA_OUT_0_4[16]\, DATA_OUT_0_4(15) => 
        \DATA_OUT_0_4[15]\, DATA_OUT_0_4(14) => 
        \DATA_OUT_0_4[14]\, DATA_OUT_0_4(13) => 
        \DATA_OUT_0_4[13]\, DATA_OUT_0_4(12) => 
        \DATA_OUT_0_4[12]\, DATA_OUT_0_4(11) => 
        \DATA_OUT_0_4[11]\, DATA_OUT_0_4(10) => 
        \DATA_OUT_0_4[10]\, DATA_OUT_0_4(9) => \DATA_OUT_0_4[9]\, 
        DATA_OUT_0_4(8) => \DATA_OUT_0_4[8]\, DATA_OUT_0_4(7) => 
        \DATA_OUT_0_4[7]\, DATA_OUT_0_4(6) => \DATA_OUT_0_4[6]\, 
        DATA_OUT_0_4(5) => \DATA_OUT_0_4[5]\, DATA_OUT_0_4(4) => 
        \DATA_OUT_0_4[4]\, DATA_OUT_0_4(3) => \DATA_OUT_0_4[3]\, 
        DATA_OUT_0_4(2) => \DATA_OUT_0_4[2]\, DATA_OUT_0_4(1) => 
        \DATA_OUT_0_4[1]\, DATA_OUT_0_4(0) => \DATA_OUT_0_4[0]\, 
        DATA_OUT_0_5(25) => \DATA_OUT_0_5[25]\, DATA_OUT_0_5(24)
         => \DATA_OUT_0_5[24]\, DATA_OUT_0_5(23) => 
        \DATA_OUT_0_5[23]\, DATA_OUT_0_5(22) => 
        \DATA_OUT_0_5[22]\, DATA_OUT_0_5(21) => 
        \DATA_OUT_0_5[21]\, DATA_OUT_0_5(20) => 
        \DATA_OUT_0_5[20]\, DATA_OUT_0_5(19) => 
        \DATA_OUT_0_5[19]\, DATA_OUT_0_5(18) => 
        \DATA_OUT_0_5[18]\, DATA_OUT_0_5(17) => 
        \DATA_OUT_0_5[17]\, DATA_OUT_0_5(16) => 
        \DATA_OUT_0_5[16]\, DATA_OUT_0_5(15) => 
        \DATA_OUT_0_5[15]\, DATA_OUT_0_5(14) => 
        \DATA_OUT_0_5[14]\, DATA_OUT_0_5(13) => 
        \DATA_OUT_0_5[13]\, DATA_OUT_0_5(12) => 
        \DATA_OUT_0_5[12]\, DATA_OUT_0_5(11) => 
        \DATA_OUT_0_5[11]\, DATA_OUT_0_5(10) => 
        \DATA_OUT_0_5[10]\, DATA_OUT_0_5(9) => \DATA_OUT_0_5[9]\, 
        DATA_OUT_0_5(8) => \DATA_OUT_0_5[8]\, DATA_OUT_0_5(7) => 
        \DATA_OUT_0_5[7]\, DATA_OUT_0_5(6) => \DATA_OUT_0_5[6]\, 
        DATA_OUT_0_5(5) => \DATA_OUT_0_5[5]\, DATA_OUT_0_5(4) => 
        \DATA_OUT_0_5[4]\, DATA_OUT_0_5(3) => \DATA_OUT_0_5[3]\, 
        DATA_OUT_0_5(2) => \DATA_OUT_0_5[2]\, DATA_OUT_0_5(1) => 
        \DATA_OUT_0_5[1]\, DATA_OUT_0_5(0) => \DATA_OUT_0_5[0]\, 
        DATA_OUT_0_6(25) => \DATA_OUT_0_6[25]\, DATA_OUT_0_6(24)
         => \DATA_OUT_0_6[24]\, DATA_OUT_0_6(23) => 
        \DATA_OUT_0_6[23]\, DATA_OUT_0_6(22) => 
        \DATA_OUT_0_6[22]\, DATA_OUT_0_6(21) => 
        \DATA_OUT_0_6[21]\, DATA_OUT_0_6(20) => 
        \DATA_OUT_0_6[20]\, DATA_OUT_0_6(19) => 
        \DATA_OUT_0_6[19]\, DATA_OUT_0_6(18) => 
        \DATA_OUT_0_6[18]\, DATA_OUT_0_6(17) => 
        \DATA_OUT_0_6[17]\, DATA_OUT_0_6(16) => 
        \DATA_OUT_0_6[16]\, DATA_OUT_0_6(15) => 
        \DATA_OUT_0_6[15]\, DATA_OUT_0_6(14) => 
        \DATA_OUT_0_6[14]\, DATA_OUT_0_6(13) => 
        \DATA_OUT_0_6[13]\, DATA_OUT_0_6(12) => 
        \DATA_OUT_0_6[12]\, DATA_OUT_0_6(11) => 
        \DATA_OUT_0_6[11]\, DATA_OUT_0_6(10) => 
        \DATA_OUT_0_6[10]\, DATA_OUT_0_6(9) => \DATA_OUT_0_6[9]\, 
        DATA_OUT_0_6(8) => \DATA_OUT_0_6[8]\, DATA_OUT_0_6(7) => 
        \DATA_OUT_0_6[7]\, DATA_OUT_0_6(6) => \DATA_OUT_0_6[6]\, 
        DATA_OUT_0_6(5) => \DATA_OUT_0_6[5]\, DATA_OUT_0_6(4) => 
        \DATA_OUT_0_6[4]\, DATA_OUT_0_6(3) => \DATA_OUT_0_6[3]\, 
        DATA_OUT_0_6(2) => \DATA_OUT_0_6[2]\, DATA_OUT_0_6(1) => 
        \DATA_OUT_0_6[1]\, DATA_OUT_0_6(0) => \DATA_OUT_0_6[0]\, 
        DATA_OUT_0_7(25) => \DATA_OUT_0_7[25]\, DATA_OUT_0_7(24)
         => \DATA_OUT_0_7[24]\, DATA_OUT_0_7(23) => 
        \DATA_OUT_0_7[23]\, DATA_OUT_0_7(22) => 
        \DATA_OUT_0_7[22]\, DATA_OUT_0_7(21) => 
        \DATA_OUT_0_7[21]\, DATA_OUT_0_7(20) => 
        \DATA_OUT_0_7[20]\, DATA_OUT_0_7(19) => 
        \DATA_OUT_0_7[19]\, DATA_OUT_0_7(18) => 
        \DATA_OUT_0_7[18]\, DATA_OUT_0_7(17) => 
        \DATA_OUT_0_7[17]\, DATA_OUT_0_7(16) => 
        \DATA_OUT_0_7[16]\, DATA_OUT_0_7(15) => 
        \DATA_OUT_0_7[15]\, DATA_OUT_0_7(14) => 
        \DATA_OUT_0_7[14]\, DATA_OUT_0_7(13) => 
        \DATA_OUT_0_7[13]\, DATA_OUT_0_7(12) => 
        \DATA_OUT_0_7[12]\, DATA_OUT_0_7(11) => 
        \DATA_OUT_0_7[11]\, DATA_OUT_0_7(10) => 
        \DATA_OUT_0_7[10]\, DATA_OUT_0_7(9) => \DATA_OUT_0_7[9]\, 
        DATA_OUT_0_7(8) => \DATA_OUT_0_7[8]\, DATA_OUT_0_7(7) => 
        \DATA_OUT_0_7[7]\, DATA_OUT_0_7(6) => \DATA_OUT_0_7[6]\, 
        DATA_OUT_0_7(5) => \DATA_OUT_0_7[5]\, DATA_OUT_0_7(4) => 
        \DATA_OUT_0_7[4]\, DATA_OUT_0_7(3) => \DATA_OUT_0_7[3]\, 
        DATA_OUT_0_7(2) => \DATA_OUT_0_7[2]\, DATA_OUT_0_7(1) => 
        \DATA_OUT_0_7[1]\, DATA_OUT_0_7(0) => \DATA_OUT_0_7[0]\, 
        DATA_OUT_0_8(25) => \DATA_OUT_0_8[25]\, DATA_OUT_0_8(24)
         => \DATA_OUT_0_8[24]\, DATA_OUT_0_8(23) => 
        \DATA_OUT_0_8[23]\, DATA_OUT_0_8(22) => 
        \DATA_OUT_0_8[22]\, DATA_OUT_0_8(21) => 
        \DATA_OUT_0_8[21]\, DATA_OUT_0_8(20) => 
        \DATA_OUT_0_8[20]\, DATA_OUT_0_8(19) => 
        \DATA_OUT_0_8[19]\, DATA_OUT_0_8(18) => 
        \DATA_OUT_0_8[18]\, DATA_OUT_0_8(17) => 
        \DATA_OUT_0_8[17]\, DATA_OUT_0_8(16) => 
        \DATA_OUT_0_8[16]\, DATA_OUT_0_8(15) => 
        \DATA_OUT_0_8[15]\, DATA_OUT_0_8(14) => 
        \DATA_OUT_0_8[14]\, DATA_OUT_0_8(13) => 
        \DATA_OUT_0_8[13]\, DATA_OUT_0_8(12) => 
        \DATA_OUT_0_8[12]\, DATA_OUT_0_8(11) => 
        \DATA_OUT_0_8[11]\, DATA_OUT_0_8(10) => 
        \DATA_OUT_0_8[10]\, DATA_OUT_0_8(9) => \DATA_OUT_0_8[9]\, 
        DATA_OUT_0_8(8) => \DATA_OUT_0_8[8]\, DATA_OUT_0_8(7) => 
        \DATA_OUT_0_8[7]\, DATA_OUT_0_8(6) => \DATA_OUT_0_8[6]\, 
        DATA_OUT_0_8(5) => \DATA_OUT_0_8[5]\, DATA_OUT_0_8(4) => 
        \DATA_OUT_0_8[4]\, DATA_OUT_0_8(3) => \DATA_OUT_0_8[3]\, 
        DATA_OUT_0_8(2) => \DATA_OUT_0_8[2]\, DATA_OUT_0_8(1) => 
        \DATA_OUT_0_8[1]\, DATA_OUT_0_8(0) => \DATA_OUT_0_8[0]\, 
        DATA_OUT_0_9(25) => \DATA_OUT_0_9[25]\, DATA_OUT_0_9(24)
         => \DATA_OUT_0_9[24]\, DATA_OUT_0_9(23) => 
        \DATA_OUT_0_9[23]\, DATA_OUT_0_9(22) => 
        \DATA_OUT_0_9[22]\, DATA_OUT_0_9(21) => 
        \DATA_OUT_0_9[21]\, DATA_OUT_0_9(20) => 
        \DATA_OUT_0_9[20]\, DATA_OUT_0_9(19) => 
        \DATA_OUT_0_9[19]\, DATA_OUT_0_9(18) => 
        \DATA_OUT_0_9[18]\, DATA_OUT_0_9(17) => 
        \DATA_OUT_0_9[17]\, DATA_OUT_0_9(16) => 
        \DATA_OUT_0_9[16]\, DATA_OUT_0_9(15) => 
        \DATA_OUT_0_9[15]\, DATA_OUT_0_9(14) => 
        \DATA_OUT_0_9[14]\, DATA_OUT_0_9(13) => 
        \DATA_OUT_0_9[13]\, DATA_OUT_0_9(12) => 
        \DATA_OUT_0_9[12]\, DATA_OUT_0_9(11) => 
        \DATA_OUT_0_9[11]\, DATA_OUT_0_9(10) => 
        \DATA_OUT_0_9[10]\, DATA_OUT_0_9(9) => \DATA_OUT_0_9[9]\, 
        DATA_OUT_0_9(8) => \DATA_OUT_0_9[8]\, DATA_OUT_0_9(7) => 
        \DATA_OUT_0_9[7]\, DATA_OUT_0_9(6) => \DATA_OUT_0_9[6]\, 
        DATA_OUT_0_9(5) => \DATA_OUT_0_9[5]\, DATA_OUT_0_9(4) => 
        \DATA_OUT_0_9[4]\, DATA_OUT_0_9(3) => \DATA_OUT_0_9[3]\, 
        DATA_OUT_0_9(2) => \DATA_OUT_0_9[2]\, DATA_OUT_0_9(1) => 
        \DATA_OUT_0_9[1]\, DATA_OUT_0_9(0) => \DATA_OUT_0_9[0]\, 
        DATA_OUT_0_26(25) => \DATA_OUT_0_26[25]\, 
        DATA_OUT_0_26(24) => \DATA_OUT_0_26[24]\, 
        DATA_OUT_0_26(23) => \DATA_OUT_0_26[23]\, 
        DATA_OUT_0_26(22) => \DATA_OUT_0_26[22]\, 
        DATA_OUT_0_26(21) => \DATA_OUT_0_26[21]\, 
        DATA_OUT_0_26(20) => \DATA_OUT_0_26[20]\, 
        DATA_OUT_0_26(19) => \DATA_OUT_0_26[19]\, 
        DATA_OUT_0_26(18) => \DATA_OUT_0_26[18]\, 
        DATA_OUT_0_26(17) => \DATA_OUT_0_26[17]\, 
        DATA_OUT_0_26(16) => \DATA_OUT_0_26[16]\, 
        DATA_OUT_0_26(15) => \DATA_OUT_0_26[15]\, 
        DATA_OUT_0_26(14) => \DATA_OUT_0_26[14]\, 
        DATA_OUT_0_26(13) => \DATA_OUT_0_26[13]\, 
        DATA_OUT_0_26(12) => \DATA_OUT_0_26[12]\, 
        DATA_OUT_0_26(11) => \DATA_OUT_0_26[11]\, 
        DATA_OUT_0_26(10) => \DATA_OUT_0_26[10]\, 
        DATA_OUT_0_26(9) => \DATA_OUT_0_26[9]\, DATA_OUT_0_26(8)
         => \DATA_OUT_0_26[8]\, DATA_OUT_0_26(7) => 
        \DATA_OUT_0_26[7]\, DATA_OUT_0_26(6) => 
        \DATA_OUT_0_26[6]\, DATA_OUT_0_26(5) => 
        \DATA_OUT_0_26[5]\, DATA_OUT_0_26(4) => 
        \DATA_OUT_0_26[4]\, DATA_OUT_0_26(3) => 
        \DATA_OUT_0_26[3]\, DATA_OUT_0_26(2) => 
        \DATA_OUT_0_26[2]\, DATA_OUT_0_26(1) => 
        \DATA_OUT_0_26[1]\, DATA_OUT_0_26(0) => 
        \DATA_OUT_0_26[0]\, DATA_OUT_0_27(25) => 
        \DATA_OUT_0_27[25]\, DATA_OUT_0_27(24) => 
        \DATA_OUT_0_27[24]\, DATA_OUT_0_27(23) => 
        \DATA_OUT_0_27[23]\, DATA_OUT_0_27(22) => 
        \DATA_OUT_0_27[22]\, DATA_OUT_0_27(21) => 
        \DATA_OUT_0_27[21]\, DATA_OUT_0_27(20) => 
        \DATA_OUT_0_27[20]\, DATA_OUT_0_27(19) => 
        \DATA_OUT_0_27[19]\, DATA_OUT_0_27(18) => 
        \DATA_OUT_0_27[18]\, DATA_OUT_0_27(17) => 
        \DATA_OUT_0_27[17]\, DATA_OUT_0_27(16) => 
        \DATA_OUT_0_27[16]\, DATA_OUT_0_27(15) => 
        \DATA_OUT_0_27[15]\, DATA_OUT_0_27(14) => 
        \DATA_OUT_0_27[14]\, DATA_OUT_0_27(13) => 
        \DATA_OUT_0_27[13]\, DATA_OUT_0_27(12) => 
        \DATA_OUT_0_27[12]\, DATA_OUT_0_27(11) => 
        \DATA_OUT_0_27[11]\, DATA_OUT_0_27(10) => 
        \DATA_OUT_0_27[10]\, DATA_OUT_0_27(9) => 
        \DATA_OUT_0_27[9]\, DATA_OUT_0_27(8) => 
        \DATA_OUT_0_27[8]\, DATA_OUT_0_27(7) => 
        \DATA_OUT_0_27[7]\, DATA_OUT_0_27(6) => 
        \DATA_OUT_0_27[6]\, DATA_OUT_0_27(5) => 
        \DATA_OUT_0_27[5]\, DATA_OUT_0_27(4) => 
        \DATA_OUT_0_27[4]\, DATA_OUT_0_27(3) => 
        \DATA_OUT_0_27[3]\, DATA_OUT_0_27(2) => 
        \DATA_OUT_0_27[2]\, DATA_OUT_0_27(1) => 
        \DATA_OUT_0_27[1]\, DATA_OUT_0_27(0) => 
        \DATA_OUT_0_27[0]\, DATA_OUT_0_28(25) => 
        \DATA_OUT_0_28[25]\, DATA_OUT_0_28(24) => 
        \DATA_OUT_0_28[24]\, DATA_OUT_0_28(23) => 
        \DATA_OUT_0_28[23]\, DATA_OUT_0_28(22) => 
        \DATA_OUT_0_28[22]\, DATA_OUT_0_28(21) => 
        \DATA_OUT_0_28[21]\, DATA_OUT_0_28(20) => 
        \DATA_OUT_0_28[20]\, DATA_OUT_0_28(19) => 
        \DATA_OUT_0_28[19]\, DATA_OUT_0_28(18) => 
        \DATA_OUT_0_28[18]\, DATA_OUT_0_28(17) => 
        \DATA_OUT_0_28[17]\, DATA_OUT_0_28(16) => 
        \DATA_OUT_0_28[16]\, DATA_OUT_0_28(15) => 
        \DATA_OUT_0_28[15]\, DATA_OUT_0_28(14) => 
        \DATA_OUT_0_28[14]\, DATA_OUT_0_28(13) => 
        \DATA_OUT_0_28[13]\, DATA_OUT_0_28(12) => 
        \DATA_OUT_0_28[12]\, DATA_OUT_0_28(11) => 
        \DATA_OUT_0_28[11]\, DATA_OUT_0_28(10) => 
        \DATA_OUT_0_28[10]\, DATA_OUT_0_28(9) => 
        \DATA_OUT_0_28[9]\, DATA_OUT_0_28(8) => 
        \DATA_OUT_0_28[8]\, DATA_OUT_0_28(7) => 
        \DATA_OUT_0_28[7]\, DATA_OUT_0_28(6) => 
        \DATA_OUT_0_28[6]\, DATA_OUT_0_28(5) => 
        \DATA_OUT_0_28[5]\, DATA_OUT_0_28(4) => 
        \DATA_OUT_0_28[4]\, DATA_OUT_0_28(3) => 
        \DATA_OUT_0_28[3]\, DATA_OUT_0_28(2) => 
        \DATA_OUT_0_28[2]\, DATA_OUT_0_28(1) => 
        \DATA_OUT_0_28[1]\, DATA_OUT_0_28(0) => 
        \DATA_OUT_0_28[0]\, DATA_OUT_0_29(25) => 
        \DATA_OUT_0_29[25]\, DATA_OUT_0_29(24) => 
        \DATA_OUT_0_29[24]\, DATA_OUT_0_29(23) => 
        \DATA_OUT_0_29[23]\, DATA_OUT_0_29(22) => 
        \DATA_OUT_0_29[22]\, DATA_OUT_0_29(21) => 
        \DATA_OUT_0_29[21]\, DATA_OUT_0_29(20) => 
        \DATA_OUT_0_29[20]\, DATA_OUT_0_29(19) => 
        \DATA_OUT_0_29[19]\, DATA_OUT_0_29(18) => 
        \DATA_OUT_0_29[18]\, DATA_OUT_0_29(17) => 
        \DATA_OUT_0_29[17]\, DATA_OUT_0_29(16) => 
        \DATA_OUT_0_29[16]\, DATA_OUT_0_29(15) => 
        \DATA_OUT_0_29[15]\, DATA_OUT_0_29(14) => 
        \DATA_OUT_0_29[14]\, DATA_OUT_0_29(13) => 
        \DATA_OUT_0_29[13]\, DATA_OUT_0_29(12) => 
        \DATA_OUT_0_29[12]\, DATA_OUT_0_29(11) => 
        \DATA_OUT_0_29[11]\, DATA_OUT_0_29(10) => 
        \DATA_OUT_0_29[10]\, DATA_OUT_0_29(9) => 
        \DATA_OUT_0_29[9]\, DATA_OUT_0_29(8) => 
        \DATA_OUT_0_29[8]\, DATA_OUT_0_29(7) => 
        \DATA_OUT_0_29[7]\, DATA_OUT_0_29(6) => 
        \DATA_OUT_0_29[6]\, DATA_OUT_0_29(5) => 
        \DATA_OUT_0_29[5]\, DATA_OUT_0_29(4) => 
        \DATA_OUT_0_29[4]\, DATA_OUT_0_29(3) => 
        \DATA_OUT_0_29[3]\, DATA_OUT_0_29(2) => 
        \DATA_OUT_0_29[2]\, DATA_OUT_0_29(1) => 
        \DATA_OUT_0_29[1]\, DATA_OUT_0_29(0) => 
        \DATA_OUT_0_29[0]\, DATA_OUT_0_30(25) => 
        \DATA_OUT_0_30[25]\, DATA_OUT_0_30(24) => 
        \DATA_OUT_0_30[24]\, DATA_OUT_0_30(23) => 
        \DATA_OUT_0_30[23]\, DATA_OUT_0_30(22) => 
        \DATA_OUT_0_30[22]\, DATA_OUT_0_30(21) => 
        \DATA_OUT_0_30[21]\, DATA_OUT_0_30(20) => 
        \DATA_OUT_0_30[20]\, DATA_OUT_0_30(19) => 
        \DATA_OUT_0_30[19]\, DATA_OUT_0_30(18) => 
        \DATA_OUT_0_30[18]\, DATA_OUT_0_30(17) => 
        \DATA_OUT_0_30[17]\, DATA_OUT_0_30(16) => 
        \DATA_OUT_0_30[16]\, DATA_OUT_0_30(15) => 
        \DATA_OUT_0_30[15]\, DATA_OUT_0_30(14) => 
        \DATA_OUT_0_30[14]\, DATA_OUT_0_30(13) => 
        \DATA_OUT_0_30[13]\, DATA_OUT_0_30(12) => 
        \DATA_OUT_0_30[12]\, DATA_OUT_0_30(11) => 
        \DATA_OUT_0_30[11]\, DATA_OUT_0_30(10) => 
        \DATA_OUT_0_30[10]\, DATA_OUT_0_30(9) => 
        \DATA_OUT_0_30[9]\, DATA_OUT_0_30(8) => 
        \DATA_OUT_0_30[8]\, DATA_OUT_0_30(7) => 
        \DATA_OUT_0_30[7]\, DATA_OUT_0_30(6) => 
        \DATA_OUT_0_30[6]\, DATA_OUT_0_30(5) => 
        \DATA_OUT_0_30[5]\, DATA_OUT_0_30(4) => 
        \DATA_OUT_0_30[4]\, DATA_OUT_0_30(3) => 
        \DATA_OUT_0_30[3]\, DATA_OUT_0_30(2) => 
        \DATA_OUT_0_30[2]\, DATA_OUT_0_30(1) => 
        \DATA_OUT_0_30[1]\, DATA_OUT_0_30(0) => 
        \DATA_OUT_0_30[0]\, DATA_OUT_0_31(25) => 
        \DATA_OUT_0_31[25]\, DATA_OUT_0_31(24) => 
        \DATA_OUT_0_31[24]\, DATA_OUT_0_31(23) => 
        \DATA_OUT_0_31[23]\, DATA_OUT_0_31(22) => 
        \DATA_OUT_0_31[22]\, DATA_OUT_0_31(21) => 
        \DATA_OUT_0_31[21]\, DATA_OUT_0_31(20) => 
        \DATA_OUT_0_31[20]\, DATA_OUT_0_31(19) => 
        \DATA_OUT_0_31[19]\, DATA_OUT_0_31(18) => 
        \DATA_OUT_0_31[18]\, DATA_OUT_0_31(17) => 
        \DATA_OUT_0_31[17]\, DATA_OUT_0_31(16) => 
        \DATA_OUT_0_31[16]\, DATA_OUT_0_31(15) => 
        \DATA_OUT_0_31[15]\, DATA_OUT_0_31(14) => 
        \DATA_OUT_0_31[14]\, DATA_OUT_0_31(13) => 
        \DATA_OUT_0_31[13]\, DATA_OUT_0_31(12) => 
        \DATA_OUT_0_31[12]\, DATA_OUT_0_31(11) => 
        \DATA_OUT_0_31[11]\, DATA_OUT_0_31(10) => 
        \DATA_OUT_0_31[10]\, DATA_OUT_0_31(9) => 
        \DATA_OUT_0_31[9]\, DATA_OUT_0_31(8) => 
        \DATA_OUT_0_31[8]\, DATA_OUT_0_31(7) => 
        \DATA_OUT_0_31[7]\, DATA_OUT_0_31(6) => 
        \DATA_OUT_0_31[6]\, DATA_OUT_0_31(5) => 
        \DATA_OUT_0_31[5]\, DATA_OUT_0_31(4) => 
        \DATA_OUT_0_31[4]\, DATA_OUT_0_31(3) => 
        \DATA_OUT_0_31[3]\, DATA_OUT_0_31(2) => 
        \DATA_OUT_0_31[2]\, DATA_OUT_0_31(1) => 
        \DATA_OUT_0_31[1]\, DATA_OUT_0_31(0) => 
        \DATA_OUT_0_31[0]\, DATA_OUT_0_32(25) => 
        \DATA_OUT_0_32[25]\, DATA_OUT_0_32(24) => 
        \DATA_OUT_0_32[24]\, DATA_OUT_0_32(23) => 
        \DATA_OUT_0_32[23]\, DATA_OUT_0_32(22) => 
        \DATA_OUT_0_32[22]\, DATA_OUT_0_32(21) => 
        \DATA_OUT_0_32[21]\, DATA_OUT_0_32(20) => 
        \DATA_OUT_0_32[20]\, DATA_OUT_0_32(19) => 
        \DATA_OUT_0_32[19]\, DATA_OUT_0_32(18) => 
        \DATA_OUT_0_32[18]\, DATA_OUT_0_32(17) => 
        \DATA_OUT_0_32[17]\, DATA_OUT_0_32(16) => 
        \DATA_OUT_0_32[16]\, DATA_OUT_0_32(15) => 
        \DATA_OUT_0_32[15]\, DATA_OUT_0_32(14) => 
        \DATA_OUT_0_32[14]\, DATA_OUT_0_32(13) => 
        \DATA_OUT_0_32[13]\, DATA_OUT_0_32(12) => 
        \DATA_OUT_0_32[12]\, DATA_OUT_0_32(11) => 
        \DATA_OUT_0_32[11]\, DATA_OUT_0_32(10) => 
        \DATA_OUT_0_32[10]\, DATA_OUT_0_32(9) => 
        \DATA_OUT_0_32[9]\, DATA_OUT_0_32(8) => 
        \DATA_OUT_0_32[8]\, DATA_OUT_0_32(7) => 
        \DATA_OUT_0_32[7]\, DATA_OUT_0_32(6) => 
        \DATA_OUT_0_32[6]\, DATA_OUT_0_32(5) => 
        \DATA_OUT_0_32[5]\, DATA_OUT_0_32(4) => 
        \DATA_OUT_0_32[4]\, DATA_OUT_0_32(3) => 
        \DATA_OUT_0_32[3]\, DATA_OUT_0_32(2) => 
        \DATA_OUT_0_32[2]\, DATA_OUT_0_32(1) => 
        \DATA_OUT_0_32[1]\, DATA_OUT_0_32(0) => 
        \DATA_OUT_0_32[0]\, DATA_OUT_0_33(25) => 
        \DATA_OUT_0_33[25]\, DATA_OUT_0_33(24) => 
        \DATA_OUT_0_33[24]\, DATA_OUT_0_33(23) => 
        \DATA_OUT_0_33[23]\, DATA_OUT_0_33(22) => 
        \DATA_OUT_0_33[22]\, DATA_OUT_0_33(21) => 
        \DATA_OUT_0_33[21]\, DATA_OUT_0_33(20) => 
        \DATA_OUT_0_33[20]\, DATA_OUT_0_33(19) => 
        \DATA_OUT_0_33[19]\, DATA_OUT_0_33(18) => 
        \DATA_OUT_0_33[18]\, DATA_OUT_0_33(17) => 
        \DATA_OUT_0_33[17]\, DATA_OUT_0_33(16) => 
        \DATA_OUT_0_33[16]\, DATA_OUT_0_33(15) => 
        \DATA_OUT_0_33[15]\, DATA_OUT_0_33(14) => 
        \DATA_OUT_0_33[14]\, DATA_OUT_0_33(13) => 
        \DATA_OUT_0_33[13]\, DATA_OUT_0_33(12) => 
        \DATA_OUT_0_33[12]\, DATA_OUT_0_33(11) => 
        \DATA_OUT_0_33[11]\, DATA_OUT_0_33(10) => 
        \DATA_OUT_0_33[10]\, DATA_OUT_0_33(9) => 
        \DATA_OUT_0_33[9]\, DATA_OUT_0_33(8) => 
        \DATA_OUT_0_33[8]\, DATA_OUT_0_33(7) => 
        \DATA_OUT_0_33[7]\, DATA_OUT_0_33(6) => 
        \DATA_OUT_0_33[6]\, DATA_OUT_0_33(5) => 
        \DATA_OUT_0_33[5]\, DATA_OUT_0_33(4) => 
        \DATA_OUT_0_33[4]\, DATA_OUT_0_33(3) => 
        \DATA_OUT_0_33[3]\, DATA_OUT_0_33(2) => 
        \DATA_OUT_0_33[2]\, DATA_OUT_0_33(1) => 
        \DATA_OUT_0_33[1]\, DATA_OUT_0_33(0) => 
        \DATA_OUT_0_33[0]\, DATA_OUT_0_34(25) => 
        \DATA_OUT_0_34[25]\, DATA_OUT_0_34(24) => 
        \DATA_OUT_0_34[24]\, DATA_OUT_0_34(23) => 
        \DATA_OUT_0_34[23]\, DATA_OUT_0_34(22) => 
        \DATA_OUT_0_34[22]\, DATA_OUT_0_34(21) => 
        \DATA_OUT_0_34[21]\, DATA_OUT_0_34(20) => 
        \DATA_OUT_0_34[20]\, DATA_OUT_0_34(19) => 
        \DATA_OUT_0_34[19]\, DATA_OUT_0_34(18) => 
        \DATA_OUT_0_34[18]\, DATA_OUT_0_34(17) => 
        \DATA_OUT_0_34[17]\, DATA_OUT_0_34(16) => 
        \DATA_OUT_0_34[16]\, DATA_OUT_0_34(15) => 
        \DATA_OUT_0_34[15]\, DATA_OUT_0_34(14) => 
        \DATA_OUT_0_34[14]\, DATA_OUT_0_34(13) => 
        \DATA_OUT_0_34[13]\, DATA_OUT_0_34(12) => 
        \DATA_OUT_0_34[12]\, DATA_OUT_0_34(11) => 
        \DATA_OUT_0_34[11]\, DATA_OUT_0_34(10) => 
        \DATA_OUT_0_34[10]\, DATA_OUT_0_34(9) => 
        \DATA_OUT_0_34[9]\, DATA_OUT_0_34(8) => 
        \DATA_OUT_0_34[8]\, DATA_OUT_0_34(7) => 
        \DATA_OUT_0_34[7]\, DATA_OUT_0_34(6) => 
        \DATA_OUT_0_34[6]\, DATA_OUT_0_34(5) => 
        \DATA_OUT_0_34[5]\, DATA_OUT_0_34(4) => 
        \DATA_OUT_0_34[4]\, DATA_OUT_0_34(3) => 
        \DATA_OUT_0_34[3]\, DATA_OUT_0_34(2) => 
        \DATA_OUT_0_34[2]\, DATA_OUT_0_34(1) => 
        \DATA_OUT_0_34[1]\, DATA_OUT_0_34(0) => 
        \DATA_OUT_0_34[0]\, DATA_OUT_0_35(25) => 
        \DATA_OUT_0_35[25]\, DATA_OUT_0_35(24) => 
        \DATA_OUT_0_35[24]\, DATA_OUT_0_35(23) => 
        \DATA_OUT_0_35[23]\, DATA_OUT_0_35(22) => 
        \DATA_OUT_0_35[22]\, DATA_OUT_0_35(21) => 
        \DATA_OUT_0_35[21]\, DATA_OUT_0_35(20) => 
        \DATA_OUT_0_35[20]\, DATA_OUT_0_35(19) => 
        \DATA_OUT_0_35[19]\, DATA_OUT_0_35(18) => 
        \DATA_OUT_0_35[18]\, DATA_OUT_0_35(17) => 
        \DATA_OUT_0_35[17]\, DATA_OUT_0_35(16) => 
        \DATA_OUT_0_35[16]\, DATA_OUT_0_35(15) => 
        \DATA_OUT_0_35[15]\, DATA_OUT_0_35(14) => 
        \DATA_OUT_0_35[14]\, DATA_OUT_0_35(13) => 
        \DATA_OUT_0_35[13]\, DATA_OUT_0_35(12) => 
        \DATA_OUT_0_35[12]\, DATA_OUT_0_35(11) => 
        \DATA_OUT_0_35[11]\, DATA_OUT_0_35(10) => 
        \DATA_OUT_0_35[10]\, DATA_OUT_0_35(9) => 
        \DATA_OUT_0_35[9]\, DATA_OUT_0_35(8) => 
        \DATA_OUT_0_35[8]\, DATA_OUT_0_35(7) => 
        \DATA_OUT_0_35[7]\, DATA_OUT_0_35(6) => 
        \DATA_OUT_0_35[6]\, DATA_OUT_0_35(5) => 
        \DATA_OUT_0_35[5]\, DATA_OUT_0_35(4) => 
        \DATA_OUT_0_35[4]\, DATA_OUT_0_35(3) => 
        \DATA_OUT_0_35[3]\, DATA_OUT_0_35(2) => 
        \DATA_OUT_0_35[2]\, DATA_OUT_0_35(1) => 
        \DATA_OUT_0_35[1]\, DATA_OUT_0_35(0) => 
        \DATA_OUT_0_35[0]\, DATA_OUT_0_36(25) => 
        \DATA_OUT_0_36[25]\, DATA_OUT_0_36(24) => 
        \DATA_OUT_0_36[24]\, DATA_OUT_0_36(23) => 
        \DATA_OUT_0_36[23]\, DATA_OUT_0_36(22) => 
        \DATA_OUT_0_36[22]\, DATA_OUT_0_36(21) => 
        \DATA_OUT_0_36[21]\, DATA_OUT_0_36(20) => 
        \DATA_OUT_0_36[20]\, DATA_OUT_0_36(19) => 
        \DATA_OUT_0_36[19]\, DATA_OUT_0_36(18) => 
        \DATA_OUT_0_36[18]\, DATA_OUT_0_36(17) => 
        \DATA_OUT_0_36[17]\, DATA_OUT_0_36(16) => 
        \DATA_OUT_0_36[16]\, DATA_OUT_0_36(15) => 
        \DATA_OUT_0_36[15]\, DATA_OUT_0_36(14) => 
        \DATA_OUT_0_36[14]\, DATA_OUT_0_36(13) => 
        \DATA_OUT_0_36[13]\, DATA_OUT_0_36(12) => 
        \DATA_OUT_0_36[12]\, DATA_OUT_0_36(11) => 
        \DATA_OUT_0_36[11]\, DATA_OUT_0_36(10) => 
        \DATA_OUT_0_36[10]\, DATA_OUT_0_36(9) => 
        \DATA_OUT_0_36[9]\, DATA_OUT_0_36(8) => 
        \DATA_OUT_0_36[8]\, DATA_OUT_0_36(7) => 
        \DATA_OUT_0_36[7]\, DATA_OUT_0_36(6) => 
        \DATA_OUT_0_36[6]\, DATA_OUT_0_36(5) => 
        \DATA_OUT_0_36[5]\, DATA_OUT_0_36(4) => 
        \DATA_OUT_0_36[4]\, DATA_OUT_0_36(3) => 
        \DATA_OUT_0_36[3]\, DATA_OUT_0_36(2) => 
        \DATA_OUT_0_36[2]\, DATA_OUT_0_36(1) => 
        \DATA_OUT_0_36[1]\, DATA_OUT_0_36(0) => 
        \DATA_OUT_0_36[0]\, DATA_OUT_0_37(25) => 
        \DATA_OUT_0_37[25]\, DATA_OUT_0_37(24) => 
        \DATA_OUT_0_37[24]\, DATA_OUT_0_37(23) => 
        \DATA_OUT_0_37[23]\, DATA_OUT_0_37(22) => 
        \DATA_OUT_0_37[22]\, DATA_OUT_0_37(21) => 
        \DATA_OUT_0_37[21]\, DATA_OUT_0_37(20) => 
        \DATA_OUT_0_37[20]\, DATA_OUT_0_37(19) => 
        \DATA_OUT_0_37[19]\, DATA_OUT_0_37(18) => 
        \DATA_OUT_0_37[18]\, DATA_OUT_0_37(17) => 
        \DATA_OUT_0_37[17]\, DATA_OUT_0_37(16) => 
        \DATA_OUT_0_37[16]\, DATA_OUT_0_37(15) => 
        \DATA_OUT_0_37[15]\, DATA_OUT_0_37(14) => 
        \DATA_OUT_0_37[14]\, DATA_OUT_0_37(13) => 
        \DATA_OUT_0_37[13]\, DATA_OUT_0_37(12) => 
        \DATA_OUT_0_37[12]\, DATA_OUT_0_37(11) => 
        \DATA_OUT_0_37[11]\, DATA_OUT_0_37(10) => 
        \DATA_OUT_0_37[10]\, DATA_OUT_0_37(9) => 
        \DATA_OUT_0_37[9]\, DATA_OUT_0_37(8) => 
        \DATA_OUT_0_37[8]\, DATA_OUT_0_37(7) => 
        \DATA_OUT_0_37[7]\, DATA_OUT_0_37(6) => 
        \DATA_OUT_0_37[6]\, DATA_OUT_0_37(5) => 
        \DATA_OUT_0_37[5]\, DATA_OUT_0_37(4) => 
        \DATA_OUT_0_37[4]\, DATA_OUT_0_37(3) => 
        \DATA_OUT_0_37[3]\, DATA_OUT_0_37(2) => 
        \DATA_OUT_0_37[2]\, DATA_OUT_0_37(1) => 
        \DATA_OUT_0_37[1]\, DATA_OUT_0_37(0) => 
        \DATA_OUT_0_37[0]\, DATA_OUT_0_38(25) => 
        \DATA_OUT_0_38[25]\, DATA_OUT_0_38(24) => 
        \DATA_OUT_0_38[24]\, DATA_OUT_0_38(23) => 
        \DATA_OUT_0_38[23]\, DATA_OUT_0_38(22) => 
        \DATA_OUT_0_38[22]\, DATA_OUT_0_38(21) => 
        \DATA_OUT_0_38[21]\, DATA_OUT_0_38(20) => 
        \DATA_OUT_0_38[20]\, DATA_OUT_0_38(19) => 
        \DATA_OUT_0_38[19]\, DATA_OUT_0_38(18) => 
        \DATA_OUT_0_38[18]\, DATA_OUT_0_38(17) => 
        \DATA_OUT_0_38[17]\, DATA_OUT_0_38(16) => 
        \DATA_OUT_0_38[16]\, DATA_OUT_0_38(15) => 
        \DATA_OUT_0_38[15]\, DATA_OUT_0_38(14) => 
        \DATA_OUT_0_38[14]\, DATA_OUT_0_38(13) => 
        \DATA_OUT_0_38[13]\, DATA_OUT_0_38(12) => 
        \DATA_OUT_0_38[12]\, DATA_OUT_0_38(11) => 
        \DATA_OUT_0_38[11]\, DATA_OUT_0_38(10) => 
        \DATA_OUT_0_38[10]\, DATA_OUT_0_38(9) => 
        \DATA_OUT_0_38[9]\, DATA_OUT_0_38(8) => 
        \DATA_OUT_0_38[8]\, DATA_OUT_0_38(7) => 
        \DATA_OUT_0_38[7]\, DATA_OUT_0_38(6) => 
        \DATA_OUT_0_38[6]\, DATA_OUT_0_38(5) => 
        \DATA_OUT_0_38[5]\, DATA_OUT_0_38(4) => 
        \DATA_OUT_0_38[4]\, DATA_OUT_0_38(3) => 
        \DATA_OUT_0_38[3]\, DATA_OUT_0_38(2) => 
        \DATA_OUT_0_38[2]\, DATA_OUT_0_38(1) => 
        \DATA_OUT_0_38[1]\, DATA_OUT_0_38(0) => 
        \DATA_OUT_0_38[0]\, DATA_OUT_0_39(25) => 
        \DATA_OUT_0_39[25]\, DATA_OUT_0_39(24) => 
        \DATA_OUT_0_39[24]\, DATA_OUT_0_39(23) => 
        \DATA_OUT_0_39[23]\, DATA_OUT_0_39(22) => 
        \DATA_OUT_0_39[22]\, DATA_OUT_0_39(21) => 
        \DATA_OUT_0_39[21]\, DATA_OUT_0_39(20) => 
        \DATA_OUT_0_39[20]\, DATA_OUT_0_39(19) => 
        \DATA_OUT_0_39[19]\, DATA_OUT_0_39(18) => 
        \DATA_OUT_0_39[18]\, DATA_OUT_0_39(17) => 
        \DATA_OUT_0_39[17]\, DATA_OUT_0_39(16) => 
        \DATA_OUT_0_39[16]\, DATA_OUT_0_39(15) => 
        \DATA_OUT_0_39[15]\, DATA_OUT_0_39(14) => 
        \DATA_OUT_0_39[14]\, DATA_OUT_0_39(13) => 
        \DATA_OUT_0_39[13]\, DATA_OUT_0_39(12) => 
        \DATA_OUT_0_39[12]\, DATA_OUT_0_39(11) => 
        \DATA_OUT_0_39[11]\, DATA_OUT_0_39(10) => 
        \DATA_OUT_0_39[10]\, DATA_OUT_0_39(9) => 
        \DATA_OUT_0_39[9]\, DATA_OUT_0_39(8) => 
        \DATA_OUT_0_39[8]\, DATA_OUT_0_39(7) => 
        \DATA_OUT_0_39[7]\, DATA_OUT_0_39(6) => 
        \DATA_OUT_0_39[6]\, DATA_OUT_0_39(5) => 
        \DATA_OUT_0_39[5]\, DATA_OUT_0_39(4) => 
        \DATA_OUT_0_39[4]\, DATA_OUT_0_39(3) => 
        \DATA_OUT_0_39[3]\, DATA_OUT_0_39(2) => 
        \DATA_OUT_0_39[2]\, DATA_OUT_0_39(1) => 
        \DATA_OUT_0_39[1]\, DATA_OUT_0_39(0) => 
        \DATA_OUT_0_39[0]\, DATA_OUT_0_40(25) => 
        \DATA_OUT_0_40[25]\, DATA_OUT_0_40(24) => 
        \DATA_OUT_0_40[24]\, DATA_OUT_0_40(23) => 
        \DATA_OUT_0_40[23]\, DATA_OUT_0_40(22) => 
        \DATA_OUT_0_40[22]\, DATA_OUT_0_40(21) => 
        \DATA_OUT_0_40[21]\, DATA_OUT_0_40(20) => 
        \DATA_OUT_0_40[20]\, DATA_OUT_0_40(19) => 
        \DATA_OUT_0_40[19]\, DATA_OUT_0_40(18) => 
        \DATA_OUT_0_40[18]\, DATA_OUT_0_40(17) => 
        \DATA_OUT_0_40[17]\, DATA_OUT_0_40(16) => 
        \DATA_OUT_0_40[16]\, DATA_OUT_0_40(15) => 
        \DATA_OUT_0_40[15]\, DATA_OUT_0_40(14) => 
        \DATA_OUT_0_40[14]\, DATA_OUT_0_40(13) => 
        \DATA_OUT_0_40[13]\, DATA_OUT_0_40(12) => 
        \DATA_OUT_0_40[12]\, DATA_OUT_0_40(11) => 
        \DATA_OUT_0_40[11]\, DATA_OUT_0_40(10) => 
        \DATA_OUT_0_40[10]\, DATA_OUT_0_40(9) => 
        \DATA_OUT_0_40[9]\, DATA_OUT_0_40(8) => 
        \DATA_OUT_0_40[8]\, DATA_OUT_0_40(7) => 
        \DATA_OUT_0_40[7]\, DATA_OUT_0_40(6) => 
        \DATA_OUT_0_40[6]\, DATA_OUT_0_40(5) => 
        \DATA_OUT_0_40[5]\, DATA_OUT_0_40(4) => 
        \DATA_OUT_0_40[4]\, DATA_OUT_0_40(3) => 
        \DATA_OUT_0_40[3]\, DATA_OUT_0_40(2) => 
        \DATA_OUT_0_40[2]\, DATA_OUT_0_40(1) => 
        \DATA_OUT_0_40[1]\, DATA_OUT_0_40(0) => 
        \DATA_OUT_0_40[0]\, DATA_OUT_0_41(25) => 
        \DATA_OUT_0_41[25]\, DATA_OUT_0_41(24) => 
        \DATA_OUT_0_41[24]\, DATA_OUT_0_41(23) => 
        \DATA_OUT_0_41[23]\, DATA_OUT_0_41(22) => 
        \DATA_OUT_0_41[22]\, DATA_OUT_0_41(21) => 
        \DATA_OUT_0_41[21]\, DATA_OUT_0_41(20) => 
        \DATA_OUT_0_41[20]\, DATA_OUT_0_41(19) => 
        \DATA_OUT_0_41[19]\, DATA_OUT_0_41(18) => 
        \DATA_OUT_0_41[18]\, DATA_OUT_0_41(17) => 
        \DATA_OUT_0_41[17]\, DATA_OUT_0_41(16) => 
        \DATA_OUT_0_41[16]\, DATA_OUT_0_41(15) => 
        \DATA_OUT_0_41[15]\, DATA_OUT_0_41(14) => 
        \DATA_OUT_0_41[14]\, DATA_OUT_0_41(13) => 
        \DATA_OUT_0_41[13]\, DATA_OUT_0_41(12) => 
        \DATA_OUT_0_41[12]\, DATA_OUT_0_41(11) => 
        \DATA_OUT_0_41[11]\, DATA_OUT_0_41(10) => 
        \DATA_OUT_0_41[10]\, DATA_OUT_0_41(9) => 
        \DATA_OUT_0_41[9]\, DATA_OUT_0_41(8) => 
        \DATA_OUT_0_41[8]\, DATA_OUT_0_41(7) => 
        \DATA_OUT_0_41[7]\, DATA_OUT_0_41(6) => 
        \DATA_OUT_0_41[6]\, DATA_OUT_0_41(5) => 
        \DATA_OUT_0_41[5]\, DATA_OUT_0_41(4) => 
        \DATA_OUT_0_41[4]\, DATA_OUT_0_41(3) => 
        \DATA_OUT_0_41[3]\, DATA_OUT_0_41(2) => 
        \DATA_OUT_0_41[2]\, DATA_OUT_0_41(1) => 
        \DATA_OUT_0_41[1]\, DATA_OUT_0_41(0) => 
        \DATA_OUT_0_41[0]\, DATA_OUT_0_42(25) => 
        \DATA_OUT_0_42[25]\, DATA_OUT_0_42(24) => 
        \DATA_OUT_0_42[24]\, DATA_OUT_0_42(23) => 
        \DATA_OUT_0_42[23]\, DATA_OUT_0_42(22) => 
        \DATA_OUT_0_42[22]\, DATA_OUT_0_42(21) => 
        \DATA_OUT_0_42[21]\, DATA_OUT_0_42(20) => 
        \DATA_OUT_0_42[20]\, DATA_OUT_0_42(19) => 
        \DATA_OUT_0_42[19]\, DATA_OUT_0_42(18) => 
        \DATA_OUT_0_42[18]\, DATA_OUT_0_42(17) => 
        \DATA_OUT_0_42[17]\, DATA_OUT_0_42(16) => 
        \DATA_OUT_0_42[16]\, DATA_OUT_0_42(15) => 
        \DATA_OUT_0_42[15]\, DATA_OUT_0_42(14) => 
        \DATA_OUT_0_42[14]\, DATA_OUT_0_42(13) => 
        \DATA_OUT_0_42[13]\, DATA_OUT_0_42(12) => 
        \DATA_OUT_0_42[12]\, DATA_OUT_0_42(11) => 
        \DATA_OUT_0_42[11]\, DATA_OUT_0_42(10) => 
        \DATA_OUT_0_42[10]\, DATA_OUT_0_42(9) => 
        \DATA_OUT_0_42[9]\, DATA_OUT_0_42(8) => 
        \DATA_OUT_0_42[8]\, DATA_OUT_0_42(7) => 
        \DATA_OUT_0_42[7]\, DATA_OUT_0_42(6) => 
        \DATA_OUT_0_42[6]\, DATA_OUT_0_42(5) => 
        \DATA_OUT_0_42[5]\, DATA_OUT_0_42(4) => 
        \DATA_OUT_0_42[4]\, DATA_OUT_0_42(3) => 
        \DATA_OUT_0_42[3]\, DATA_OUT_0_42(2) => 
        \DATA_OUT_0_42[2]\, DATA_OUT_0_42(1) => 
        \DATA_OUT_0_42[1]\, DATA_OUT_0_42(0) => 
        \DATA_OUT_0_42[0]\, DATA_OUT_0_43(25) => 
        \DATA_OUT_0_43[25]\, DATA_OUT_0_43(24) => 
        \DATA_OUT_0_43[24]\, DATA_OUT_0_43(23) => 
        \DATA_OUT_0_43[23]\, DATA_OUT_0_43(22) => 
        \DATA_OUT_0_43[22]\, DATA_OUT_0_43(21) => 
        \DATA_OUT_0_43[21]\, DATA_OUT_0_43(20) => 
        \DATA_OUT_0_43[20]\, DATA_OUT_0_43(19) => 
        \DATA_OUT_0_43[19]\, DATA_OUT_0_43(18) => 
        \DATA_OUT_0_43[18]\, DATA_OUT_0_43(17) => 
        \DATA_OUT_0_43[17]\, DATA_OUT_0_43(16) => 
        \DATA_OUT_0_43[16]\, DATA_OUT_0_43(15) => 
        \DATA_OUT_0_43[15]\, DATA_OUT_0_43(14) => 
        \DATA_OUT_0_43[14]\, DATA_OUT_0_43(13) => 
        \DATA_OUT_0_43[13]\, DATA_OUT_0_43(12) => 
        \DATA_OUT_0_43[12]\, DATA_OUT_0_43(11) => 
        \DATA_OUT_0_43[11]\, DATA_OUT_0_43(10) => 
        \DATA_OUT_0_43[10]\, DATA_OUT_0_43(9) => 
        \DATA_OUT_0_43[9]\, DATA_OUT_0_43(8) => 
        \DATA_OUT_0_43[8]\, DATA_OUT_0_43(7) => 
        \DATA_OUT_0_43[7]\, DATA_OUT_0_43(6) => 
        \DATA_OUT_0_43[6]\, DATA_OUT_0_43(5) => 
        \DATA_OUT_0_43[5]\, DATA_OUT_0_43(4) => 
        \DATA_OUT_0_43[4]\, DATA_OUT_0_43(3) => 
        \DATA_OUT_0_43[3]\, DATA_OUT_0_43(2) => 
        \DATA_OUT_0_43[2]\, DATA_OUT_0_43(1) => 
        \DATA_OUT_0_43[1]\, DATA_OUT_0_43(0) => 
        \DATA_OUT_0_43[0]\, DATA_OUT_0_44(25) => 
        \DATA_OUT_0_44[25]\, DATA_OUT_0_44(24) => 
        \DATA_OUT_0_44[24]\, DATA_OUT_0_44(23) => 
        \DATA_OUT_0_44[23]\, DATA_OUT_0_44(22) => 
        \DATA_OUT_0_44[22]\, DATA_OUT_0_44(21) => 
        \DATA_OUT_0_44[21]\, DATA_OUT_0_44(20) => 
        \DATA_OUT_0_44[20]\, DATA_OUT_0_44(19) => 
        \DATA_OUT_0_44[19]\, DATA_OUT_0_44(18) => 
        \DATA_OUT_0_44[18]\, DATA_OUT_0_44(17) => 
        \DATA_OUT_0_44[17]\, DATA_OUT_0_44(16) => 
        \DATA_OUT_0_44[16]\, DATA_OUT_0_44(15) => 
        \DATA_OUT_0_44[15]\, DATA_OUT_0_44(14) => 
        \DATA_OUT_0_44[14]\, DATA_OUT_0_44(13) => 
        \DATA_OUT_0_44[13]\, DATA_OUT_0_44(12) => 
        \DATA_OUT_0_44[12]\, DATA_OUT_0_44(11) => 
        \DATA_OUT_0_44[11]\, DATA_OUT_0_44(10) => 
        \DATA_OUT_0_44[10]\, DATA_OUT_0_44(9) => 
        \DATA_OUT_0_44[9]\, DATA_OUT_0_44(8) => 
        \DATA_OUT_0_44[8]\, DATA_OUT_0_44(7) => 
        \DATA_OUT_0_44[7]\, DATA_OUT_0_44(6) => 
        \DATA_OUT_0_44[6]\, DATA_OUT_0_44(5) => 
        \DATA_OUT_0_44[5]\, DATA_OUT_0_44(4) => 
        \DATA_OUT_0_44[4]\, DATA_OUT_0_44(3) => 
        \DATA_OUT_0_44[3]\, DATA_OUT_0_44(2) => 
        \DATA_OUT_0_44[2]\, DATA_OUT_0_44(1) => 
        \DATA_OUT_0_44[1]\, DATA_OUT_0_44(0) => 
        \DATA_OUT_0_44[0]\, DATA_OUT_0_45(25) => 
        \DATA_OUT_0_45[25]\, DATA_OUT_0_45(24) => 
        \DATA_OUT_0_45[24]\, DATA_OUT_0_45(23) => 
        \DATA_OUT_0_45[23]\, DATA_OUT_0_45(22) => 
        \DATA_OUT_0_45[22]\, DATA_OUT_0_45(21) => 
        \DATA_OUT_0_45[21]\, DATA_OUT_0_45(20) => 
        \DATA_OUT_0_45[20]\, DATA_OUT_0_45(19) => 
        \DATA_OUT_0_45[19]\, DATA_OUT_0_45(18) => 
        \DATA_OUT_0_45[18]\, DATA_OUT_0_45(17) => 
        \DATA_OUT_0_45[17]\, DATA_OUT_0_45(16) => 
        \DATA_OUT_0_45[16]\, DATA_OUT_0_45(15) => 
        \DATA_OUT_0_45[15]\, DATA_OUT_0_45(14) => 
        \DATA_OUT_0_45[14]\, DATA_OUT_0_45(13) => 
        \DATA_OUT_0_45[13]\, DATA_OUT_0_45(12) => 
        \DATA_OUT_0_45[12]\, DATA_OUT_0_45(11) => 
        \DATA_OUT_0_45[11]\, DATA_OUT_0_45(10) => 
        \DATA_OUT_0_45[10]\, DATA_OUT_0_45(9) => 
        \DATA_OUT_0_45[9]\, DATA_OUT_0_45(8) => 
        \DATA_OUT_0_45[8]\, DATA_OUT_0_45(7) => 
        \DATA_OUT_0_45[7]\, DATA_OUT_0_45(6) => 
        \DATA_OUT_0_45[6]\, DATA_OUT_0_45(5) => 
        \DATA_OUT_0_45[5]\, DATA_OUT_0_45(4) => 
        \DATA_OUT_0_45[4]\, DATA_OUT_0_45(3) => 
        \DATA_OUT_0_45[3]\, DATA_OUT_0_45(2) => 
        \DATA_OUT_0_45[2]\, DATA_OUT_0_45(1) => 
        \DATA_OUT_0_45[1]\, DATA_OUT_0_45(0) => 
        \DATA_OUT_0_45[0]\, DATA_OUT_0_46(25) => 
        \DATA_OUT_0_46[25]\, DATA_OUT_0_46(24) => 
        \DATA_OUT_0_46[24]\, DATA_OUT_0_46(23) => 
        \DATA_OUT_0_46[23]\, DATA_OUT_0_46(22) => 
        \DATA_OUT_0_46[22]\, DATA_OUT_0_46(21) => 
        \DATA_OUT_0_46[21]\, DATA_OUT_0_46(20) => 
        \DATA_OUT_0_46[20]\, DATA_OUT_0_46(19) => 
        \DATA_OUT_0_46[19]\, DATA_OUT_0_46(18) => 
        \DATA_OUT_0_46[18]\, DATA_OUT_0_46(17) => 
        \DATA_OUT_0_46[17]\, DATA_OUT_0_46(16) => 
        \DATA_OUT_0_46[16]\, DATA_OUT_0_46(15) => 
        \DATA_OUT_0_46[15]\, DATA_OUT_0_46(14) => 
        \DATA_OUT_0_46[14]\, DATA_OUT_0_46(13) => 
        \DATA_OUT_0_46[13]\, DATA_OUT_0_46(12) => 
        \DATA_OUT_0_46[12]\, DATA_OUT_0_46(11) => 
        \DATA_OUT_0_46[11]\, DATA_OUT_0_46(10) => 
        \DATA_OUT_0_46[10]\, DATA_OUT_0_46(9) => 
        \DATA_OUT_0_46[9]\, DATA_OUT_0_46(8) => 
        \DATA_OUT_0_46[8]\, DATA_OUT_0_46(7) => 
        \DATA_OUT_0_46[7]\, DATA_OUT_0_46(6) => 
        \DATA_OUT_0_46[6]\, DATA_OUT_0_46(5) => 
        \DATA_OUT_0_46[5]\, DATA_OUT_0_46(4) => 
        \DATA_OUT_0_46[4]\, DATA_OUT_0_46(3) => 
        \DATA_OUT_0_46[3]\, DATA_OUT_0_46(2) => 
        \DATA_OUT_0_46[2]\, DATA_OUT_0_46(1) => 
        \DATA_OUT_0_46[1]\, DATA_OUT_0_46(0) => 
        \DATA_OUT_0_46[0]\, DATA_OUT_0_47(25) => 
        \DATA_OUT_0_47[25]\, DATA_OUT_0_47(24) => 
        \DATA_OUT_0_47[24]\, DATA_OUT_0_47(23) => 
        \DATA_OUT_0_47[23]\, DATA_OUT_0_47(22) => 
        \DATA_OUT_0_47[22]\, DATA_OUT_0_47(21) => 
        \DATA_OUT_0_47[21]\, DATA_OUT_0_47(20) => 
        \DATA_OUT_0_47[20]\, DATA_OUT_0_47(19) => 
        \DATA_OUT_0_47[19]\, DATA_OUT_0_47(18) => 
        \DATA_OUT_0_47[18]\, DATA_OUT_0_47(17) => 
        \DATA_OUT_0_47[17]\, DATA_OUT_0_47(16) => 
        \DATA_OUT_0_47[16]\, DATA_OUT_0_47(15) => 
        \DATA_OUT_0_47[15]\, DATA_OUT_0_47(14) => 
        \DATA_OUT_0_47[14]\, DATA_OUT_0_47(13) => 
        \DATA_OUT_0_47[13]\, DATA_OUT_0_47(12) => 
        \DATA_OUT_0_47[12]\, DATA_OUT_0_47(11) => 
        \DATA_OUT_0_47[11]\, DATA_OUT_0_47(10) => 
        \DATA_OUT_0_47[10]\, DATA_OUT_0_47(9) => 
        \DATA_OUT_0_47[9]\, DATA_OUT_0_47(8) => 
        \DATA_OUT_0_47[8]\, DATA_OUT_0_47(7) => 
        \DATA_OUT_0_47[7]\, DATA_OUT_0_47(6) => 
        \DATA_OUT_0_47[6]\, DATA_OUT_0_47(5) => 
        \DATA_OUT_0_47[5]\, DATA_OUT_0_47(4) => 
        \DATA_OUT_0_47[4]\, DATA_OUT_0_47(3) => 
        \DATA_OUT_0_47[3]\, DATA_OUT_0_47(2) => 
        \DATA_OUT_0_47[2]\, DATA_OUT_0_47(1) => 
        \DATA_OUT_0_47[1]\, DATA_OUT_0_47(0) => 
        \DATA_OUT_0_47[0]\, DATA_OUT_0_48(25) => 
        \DATA_OUT_0_48[25]\, DATA_OUT_0_48(24) => 
        \DATA_OUT_0_48[24]\, DATA_OUT_0_48(23) => 
        \DATA_OUT_0_48[23]\, DATA_OUT_0_48(22) => 
        \DATA_OUT_0_48[22]\, DATA_OUT_0_48(21) => 
        \DATA_OUT_0_48[21]\, DATA_OUT_0_48(20) => 
        \DATA_OUT_0_48[20]\, DATA_OUT_0_48(19) => 
        \DATA_OUT_0_48[19]\, DATA_OUT_0_48(18) => 
        \DATA_OUT_0_48[18]\, DATA_OUT_0_48(17) => 
        \DATA_OUT_0_48[17]\, DATA_OUT_0_48(16) => 
        \DATA_OUT_0_48[16]\, DATA_OUT_0_48(15) => 
        \DATA_OUT_0_48[15]\, DATA_OUT_0_48(14) => 
        \DATA_OUT_0_48[14]\, DATA_OUT_0_48(13) => 
        \DATA_OUT_0_48[13]\, DATA_OUT_0_48(12) => 
        \DATA_OUT_0_48[12]\, DATA_OUT_0_48(11) => 
        \DATA_OUT_0_48[11]\, DATA_OUT_0_48(10) => 
        \DATA_OUT_0_48[10]\, DATA_OUT_0_48(9) => 
        \DATA_OUT_0_48[9]\, DATA_OUT_0_48(8) => 
        \DATA_OUT_0_48[8]\, DATA_OUT_0_48(7) => 
        \DATA_OUT_0_48[7]\, DATA_OUT_0_48(6) => 
        \DATA_OUT_0_48[6]\, DATA_OUT_0_48(5) => 
        \DATA_OUT_0_48[5]\, DATA_OUT_0_48(4) => 
        \DATA_OUT_0_48[4]\, DATA_OUT_0_48(3) => 
        \DATA_OUT_0_48[3]\, DATA_OUT_0_48(2) => 
        \DATA_OUT_0_48[2]\, DATA_OUT_0_48(1) => 
        \DATA_OUT_0_48[1]\, DATA_OUT_0_48(0) => 
        \DATA_OUT_0_48[0]\, DATA_OUT_0_49(25) => 
        \DATA_OUT_0_49[25]\, DATA_OUT_0_49(24) => 
        \DATA_OUT_0_49[24]\, DATA_OUT_0_49(23) => 
        \DATA_OUT_0_49[23]\, DATA_OUT_0_49(22) => 
        \DATA_OUT_0_49[22]\, DATA_OUT_0_49(21) => 
        \DATA_OUT_0_49[21]\, DATA_OUT_0_49(20) => 
        \DATA_OUT_0_49[20]\, DATA_OUT_0_49(19) => 
        \DATA_OUT_0_49[19]\, DATA_OUT_0_49(18) => 
        \DATA_OUT_0_49[18]\, DATA_OUT_0_49(17) => 
        \DATA_OUT_0_49[17]\, DATA_OUT_0_49(16) => 
        \DATA_OUT_0_49[16]\, DATA_OUT_0_49(15) => 
        \DATA_OUT_0_49[15]\, DATA_OUT_0_49(14) => 
        \DATA_OUT_0_49[14]\, DATA_OUT_0_49(13) => 
        \DATA_OUT_0_49[13]\, DATA_OUT_0_49(12) => 
        \DATA_OUT_0_49[12]\, DATA_OUT_0_49(11) => 
        \DATA_OUT_0_49[11]\, DATA_OUT_0_49(10) => 
        \DATA_OUT_0_49[10]\, DATA_OUT_0_49(9) => 
        \DATA_OUT_0_49[9]\, DATA_OUT_0_49(8) => 
        \DATA_OUT_0_49[8]\, DATA_OUT_0_49(7) => 
        \DATA_OUT_0_49[7]\, DATA_OUT_0_49(6) => 
        \DATA_OUT_0_49[6]\, DATA_OUT_0_49(5) => 
        \DATA_OUT_0_49[5]\, DATA_OUT_0_49(4) => 
        \DATA_OUT_0_49[4]\, DATA_OUT_0_49(3) => 
        \DATA_OUT_0_49[3]\, DATA_OUT_0_49(2) => 
        \DATA_OUT_0_49[2]\, DATA_OUT_0_49(1) => 
        \DATA_OUT_0_49[1]\, DATA_OUT_0_49(0) => 
        \DATA_OUT_0_49[0]\, DATA_OUT_0_50(25) => 
        \DATA_OUT_0_50[25]\, DATA_OUT_0_50(24) => 
        \DATA_OUT_0_50[24]\, DATA_OUT_0_50(23) => 
        \DATA_OUT_0_50[23]\, DATA_OUT_0_50(22) => 
        \DATA_OUT_0_50[22]\, DATA_OUT_0_50(21) => 
        \DATA_OUT_0_50[21]\, DATA_OUT_0_50(20) => 
        \DATA_OUT_0_50[20]\, DATA_OUT_0_50(19) => 
        \DATA_OUT_0_50[19]\, DATA_OUT_0_50(18) => 
        \DATA_OUT_0_50[18]\, DATA_OUT_0_50(17) => 
        \DATA_OUT_0_50[17]\, DATA_OUT_0_50(16) => 
        \DATA_OUT_0_50[16]\, DATA_OUT_0_50(15) => 
        \DATA_OUT_0_50[15]\, DATA_OUT_0_50(14) => 
        \DATA_OUT_0_50[14]\, DATA_OUT_0_50(13) => 
        \DATA_OUT_0_50[13]\, DATA_OUT_0_50(12) => 
        \DATA_OUT_0_50[12]\, DATA_OUT_0_50(11) => 
        \DATA_OUT_0_50[11]\, DATA_OUT_0_50(10) => 
        \DATA_OUT_0_50[10]\, DATA_OUT_0_50(9) => 
        \DATA_OUT_0_50[9]\, DATA_OUT_0_50(8) => 
        \DATA_OUT_0_50[8]\, DATA_OUT_0_50(7) => 
        \DATA_OUT_0_50[7]\, DATA_OUT_0_50(6) => 
        \DATA_OUT_0_50[6]\, DATA_OUT_0_50(5) => 
        \DATA_OUT_0_50[5]\, DATA_OUT_0_50(4) => 
        \DATA_OUT_0_50[4]\, DATA_OUT_0_50(3) => 
        \DATA_OUT_0_50[3]\, DATA_OUT_0_50(2) => 
        \DATA_OUT_0_50[2]\, DATA_OUT_0_50(1) => 
        \DATA_OUT_0_50[1]\, DATA_OUT_0_50(0) => 
        \DATA_OUT_0_50[0]\, DATA_OUT_0_51(25) => 
        \DATA_OUT_0_51[25]\, DATA_OUT_0_51(24) => 
        \DATA_OUT_0_51[24]\, DATA_OUT_0_51(23) => 
        \DATA_OUT_0_51[23]\, DATA_OUT_0_51(22) => 
        \DATA_OUT_0_51[22]\, DATA_OUT_0_51(21) => 
        \DATA_OUT_0_51[21]\, DATA_OUT_0_51(20) => 
        \DATA_OUT_0_51[20]\, DATA_OUT_0_51(19) => 
        \DATA_OUT_0_51[19]\, DATA_OUT_0_51(18) => 
        \DATA_OUT_0_51[18]\, DATA_OUT_0_51(17) => 
        \DATA_OUT_0_51[17]\, DATA_OUT_0_51(16) => 
        \DATA_OUT_0_51[16]\, DATA_OUT_0_51(15) => 
        \DATA_OUT_0_51[15]\, DATA_OUT_0_51(14) => 
        \DATA_OUT_0_51[14]\, DATA_OUT_0_51(13) => 
        \DATA_OUT_0_51[13]\, DATA_OUT_0_51(12) => 
        \DATA_OUT_0_51[12]\, DATA_OUT_0_51(11) => 
        \DATA_OUT_0_51[11]\, DATA_OUT_0_51(10) => 
        \DATA_OUT_0_51[10]\, DATA_OUT_0_51(9) => 
        \DATA_OUT_0_51[9]\, DATA_OUT_0_51(8) => 
        \DATA_OUT_0_51[8]\, DATA_OUT_0_51(7) => 
        \DATA_OUT_0_51[7]\, DATA_OUT_0_51(6) => 
        \DATA_OUT_0_51[6]\, DATA_OUT_0_51(5) => 
        \DATA_OUT_0_51[5]\, DATA_OUT_0_51(4) => 
        \DATA_OUT_0_51[4]\, DATA_OUT_0_51(3) => 
        \DATA_OUT_0_51[3]\, DATA_OUT_0_51(2) => 
        \DATA_OUT_0_51[2]\, DATA_OUT_0_51(1) => 
        \DATA_OUT_0_51[1]\, DATA_OUT_0_51(0) => 
        \DATA_OUT_0_51[0]\, DATA_OUT_1_0(25) => 
        \DATA_OUT_1_0[25]\, DATA_OUT_1_0(24) => 
        \DATA_OUT_1_0[24]\, DATA_OUT_1_0(23) => 
        \DATA_OUT_1_0[23]\, DATA_OUT_1_0(22) => 
        \DATA_OUT_1_0[22]\, DATA_OUT_1_0(21) => 
        \DATA_OUT_1_0[21]\, DATA_OUT_1_0(20) => 
        \DATA_OUT_1_0[20]\, DATA_OUT_1_0(19) => 
        \DATA_OUT_1_0[19]\, DATA_OUT_1_0(18) => 
        \DATA_OUT_1_0[18]\, DATA_OUT_1_0(17) => 
        \DATA_OUT_1_0[17]\, DATA_OUT_1_0(16) => 
        \DATA_OUT_1_0[16]\, DATA_OUT_1_0(15) => 
        \DATA_OUT_1_0[15]\, DATA_OUT_1_0(14) => 
        \DATA_OUT_1_0[14]\, DATA_OUT_1_0(13) => 
        \DATA_OUT_1_0[13]\, DATA_OUT_1_0(12) => 
        \DATA_OUT_1_0[12]\, DATA_OUT_1_0(11) => 
        \DATA_OUT_1_0[11]\, DATA_OUT_1_0(10) => 
        \DATA_OUT_1_0[10]\, DATA_OUT_1_0(9) => \DATA_OUT_1_0[9]\, 
        DATA_OUT_1_0(8) => \DATA_OUT_1_0[8]\, DATA_OUT_1_0(7) => 
        \DATA_OUT_1_0[7]\, DATA_OUT_1_0(6) => \DATA_OUT_1_0[6]\, 
        DATA_OUT_1_0(5) => \DATA_OUT_1_0[5]\, DATA_OUT_1_0(4) => 
        \DATA_OUT_1_0[4]\, DATA_OUT_1_0(3) => \DATA_OUT_1_0[3]\, 
        DATA_OUT_1_0(2) => \DATA_OUT_1_0[2]\, DATA_OUT_1_0(1) => 
        \DATA_OUT_1_0[1]\, DATA_OUT_1_0(0) => \DATA_OUT_1_0[0]\, 
        DATA_OUT_1_1(25) => \DATA_OUT_1_1[25]\, DATA_OUT_1_1(24)
         => \DATA_OUT_1_1[24]\, DATA_OUT_1_1(23) => 
        \DATA_OUT_1_1[23]\, DATA_OUT_1_1(22) => 
        \DATA_OUT_1_1[22]\, DATA_OUT_1_1(21) => 
        \DATA_OUT_1_1[21]\, DATA_OUT_1_1(20) => 
        \DATA_OUT_1_1[20]\, DATA_OUT_1_1(19) => 
        \DATA_OUT_1_1[19]\, DATA_OUT_1_1(18) => 
        \DATA_OUT_1_1[18]\, DATA_OUT_1_1(17) => 
        \DATA_OUT_1_1[17]\, DATA_OUT_1_1(16) => 
        \DATA_OUT_1_1[16]\, DATA_OUT_1_1(15) => 
        \DATA_OUT_1_1[15]\, DATA_OUT_1_1(14) => 
        \DATA_OUT_1_1[14]\, DATA_OUT_1_1(13) => 
        \DATA_OUT_1_1[13]\, DATA_OUT_1_1(12) => 
        \DATA_OUT_1_1[12]\, DATA_OUT_1_1(11) => 
        \DATA_OUT_1_1[11]\, DATA_OUT_1_1(10) => 
        \DATA_OUT_1_1[10]\, DATA_OUT_1_1(9) => \DATA_OUT_1_1[9]\, 
        DATA_OUT_1_1(8) => \DATA_OUT_1_1[8]\, DATA_OUT_1_1(7) => 
        \DATA_OUT_1_1[7]\, DATA_OUT_1_1(6) => \DATA_OUT_1_1[6]\, 
        DATA_OUT_1_1(5) => \DATA_OUT_1_1[5]\, DATA_OUT_1_1(4) => 
        \DATA_OUT_1_1[4]\, DATA_OUT_1_1(3) => \DATA_OUT_1_1[3]\, 
        DATA_OUT_1_1(2) => \DATA_OUT_1_1[2]\, DATA_OUT_1_1(1) => 
        \DATA_OUT_1_1[1]\, DATA_OUT_1_1(0) => \DATA_OUT_1_1[0]\, 
        DATA_OUT_1_2(25) => \DATA_OUT_1_2[25]\, DATA_OUT_1_2(24)
         => \DATA_OUT_1_2[24]\, DATA_OUT_1_2(23) => 
        \DATA_OUT_1_2[23]\, DATA_OUT_1_2(22) => 
        \DATA_OUT_1_2[22]\, DATA_OUT_1_2(21) => 
        \DATA_OUT_1_2[21]\, DATA_OUT_1_2(20) => 
        \DATA_OUT_1_2[20]\, DATA_OUT_1_2(19) => 
        \DATA_OUT_1_2[19]\, DATA_OUT_1_2(18) => 
        \DATA_OUT_1_2[18]\, DATA_OUT_1_2(17) => 
        \DATA_OUT_1_2[17]\, DATA_OUT_1_2(16) => 
        \DATA_OUT_1_2[16]\, DATA_OUT_1_2(15) => 
        \DATA_OUT_1_2[15]\, DATA_OUT_1_2(14) => 
        \DATA_OUT_1_2[14]\, DATA_OUT_1_2(13) => 
        \DATA_OUT_1_2[13]\, DATA_OUT_1_2(12) => 
        \DATA_OUT_1_2[12]\, DATA_OUT_1_2(11) => 
        \DATA_OUT_1_2[11]\, DATA_OUT_1_2(10) => 
        \DATA_OUT_1_2[10]\, DATA_OUT_1_2(9) => \DATA_OUT_1_2[9]\, 
        DATA_OUT_1_2(8) => \DATA_OUT_1_2[8]\, DATA_OUT_1_2(7) => 
        \DATA_OUT_1_2[7]\, DATA_OUT_1_2(6) => \DATA_OUT_1_2[6]\, 
        DATA_OUT_1_2(5) => \DATA_OUT_1_2[5]\, DATA_OUT_1_2(4) => 
        \DATA_OUT_1_2[4]\, DATA_OUT_1_2(3) => \DATA_OUT_1_2[3]\, 
        DATA_OUT_1_2(2) => \DATA_OUT_1_2[2]\, DATA_OUT_1_2(1) => 
        \DATA_OUT_1_2[1]\, DATA_OUT_1_2(0) => \DATA_OUT_1_2[0]\, 
        DATA_OUT_1_3(25) => \DATA_OUT_1_3[25]\, DATA_OUT_1_3(24)
         => \DATA_OUT_1_3[24]\, DATA_OUT_1_3(23) => 
        \DATA_OUT_1_3[23]\, DATA_OUT_1_3(22) => 
        \DATA_OUT_1_3[22]\, DATA_OUT_1_3(21) => 
        \DATA_OUT_1_3[21]\, DATA_OUT_1_3(20) => 
        \DATA_OUT_1_3[20]\, DATA_OUT_1_3(19) => 
        \DATA_OUT_1_3[19]\, DATA_OUT_1_3(18) => 
        \DATA_OUT_1_3[18]\, DATA_OUT_1_3(17) => 
        \DATA_OUT_1_3[17]\, DATA_OUT_1_3(16) => 
        \DATA_OUT_1_3[16]\, DATA_OUT_1_3(15) => 
        \DATA_OUT_1_3[15]\, DATA_OUT_1_3(14) => 
        \DATA_OUT_1_3[14]\, DATA_OUT_1_3(13) => 
        \DATA_OUT_1_3[13]\, DATA_OUT_1_3(12) => 
        \DATA_OUT_1_3[12]\, DATA_OUT_1_3(11) => 
        \DATA_OUT_1_3[11]\, DATA_OUT_1_3(10) => 
        \DATA_OUT_1_3[10]\, DATA_OUT_1_3(9) => \DATA_OUT_1_3[9]\, 
        DATA_OUT_1_3(8) => \DATA_OUT_1_3[8]\, DATA_OUT_1_3(7) => 
        \DATA_OUT_1_3[7]\, DATA_OUT_1_3(6) => \DATA_OUT_1_3[6]\, 
        DATA_OUT_1_3(5) => \DATA_OUT_1_3[5]\, DATA_OUT_1_3(4) => 
        \DATA_OUT_1_3[4]\, DATA_OUT_1_3(3) => \DATA_OUT_1_3[3]\, 
        DATA_OUT_1_3(2) => \DATA_OUT_1_3[2]\, DATA_OUT_1_3(1) => 
        \DATA_OUT_1_3[1]\, DATA_OUT_1_3(0) => \DATA_OUT_1_3[0]\, 
        DATA_OUT_1_4(25) => \DATA_OUT_1_4[25]\, DATA_OUT_1_4(24)
         => \DATA_OUT_1_4[24]\, DATA_OUT_1_4(23) => 
        \DATA_OUT_1_4[23]\, DATA_OUT_1_4(22) => 
        \DATA_OUT_1_4[22]\, DATA_OUT_1_4(21) => 
        \DATA_OUT_1_4[21]\, DATA_OUT_1_4(20) => 
        \DATA_OUT_1_4[20]\, DATA_OUT_1_4(19) => 
        \DATA_OUT_1_4[19]\, DATA_OUT_1_4(18) => 
        \DATA_OUT_1_4[18]\, DATA_OUT_1_4(17) => 
        \DATA_OUT_1_4[17]\, DATA_OUT_1_4(16) => 
        \DATA_OUT_1_4[16]\, DATA_OUT_1_4(15) => 
        \DATA_OUT_1_4[15]\, DATA_OUT_1_4(14) => 
        \DATA_OUT_1_4[14]\, DATA_OUT_1_4(13) => 
        \DATA_OUT_1_4[13]\, DATA_OUT_1_4(12) => 
        \DATA_OUT_1_4[12]\, DATA_OUT_1_4(11) => 
        \DATA_OUT_1_4[11]\, DATA_OUT_1_4(10) => 
        \DATA_OUT_1_4[10]\, DATA_OUT_1_4(9) => \DATA_OUT_1_4[9]\, 
        DATA_OUT_1_4(8) => \DATA_OUT_1_4[8]\, DATA_OUT_1_4(7) => 
        \DATA_OUT_1_4[7]\, DATA_OUT_1_4(6) => \DATA_OUT_1_4[6]\, 
        DATA_OUT_1_4(5) => \DATA_OUT_1_4[5]\, DATA_OUT_1_4(4) => 
        \DATA_OUT_1_4[4]\, DATA_OUT_1_4(3) => \DATA_OUT_1_4[3]\, 
        DATA_OUT_1_4(2) => \DATA_OUT_1_4[2]\, DATA_OUT_1_4(1) => 
        \DATA_OUT_1_4[1]\, DATA_OUT_1_4(0) => \DATA_OUT_1_4[0]\, 
        DATA_OUT_1_5(25) => \DATA_OUT_1_5[25]\, DATA_OUT_1_5(24)
         => \DATA_OUT_1_5[24]\, DATA_OUT_1_5(23) => 
        \DATA_OUT_1_5[23]\, DATA_OUT_1_5(22) => 
        \DATA_OUT_1_5[22]\, DATA_OUT_1_5(21) => 
        \DATA_OUT_1_5[21]\, DATA_OUT_1_5(20) => 
        \DATA_OUT_1_5[20]\, DATA_OUT_1_5(19) => 
        \DATA_OUT_1_5[19]\, DATA_OUT_1_5(18) => 
        \DATA_OUT_1_5[18]\, DATA_OUT_1_5(17) => 
        \DATA_OUT_1_5[17]\, DATA_OUT_1_5(16) => 
        \DATA_OUT_1_5[16]\, DATA_OUT_1_5(15) => 
        \DATA_OUT_1_5[15]\, DATA_OUT_1_5(14) => 
        \DATA_OUT_1_5[14]\, DATA_OUT_1_5(13) => 
        \DATA_OUT_1_5[13]\, DATA_OUT_1_5(12) => 
        \DATA_OUT_1_5[12]\, DATA_OUT_1_5(11) => 
        \DATA_OUT_1_5[11]\, DATA_OUT_1_5(10) => 
        \DATA_OUT_1_5[10]\, DATA_OUT_1_5(9) => \DATA_OUT_1_5[9]\, 
        DATA_OUT_1_5(8) => \DATA_OUT_1_5[8]\, DATA_OUT_1_5(7) => 
        \DATA_OUT_1_5[7]\, DATA_OUT_1_5(6) => \DATA_OUT_1_5[6]\, 
        DATA_OUT_1_5(5) => \DATA_OUT_1_5[5]\, DATA_OUT_1_5(4) => 
        \DATA_OUT_1_5[4]\, DATA_OUT_1_5(3) => \DATA_OUT_1_5[3]\, 
        DATA_OUT_1_5(2) => \DATA_OUT_1_5[2]\, DATA_OUT_1_5(1) => 
        \DATA_OUT_1_5[1]\, DATA_OUT_1_5(0) => \DATA_OUT_1_5[0]\, 
        DATA_OUT_1_6(25) => \DATA_OUT_1_6[25]\, DATA_OUT_1_6(24)
         => \DATA_OUT_1_6[24]\, DATA_OUT_1_6(23) => 
        \DATA_OUT_1_6[23]\, DATA_OUT_1_6(22) => 
        \DATA_OUT_1_6[22]\, DATA_OUT_1_6(21) => 
        \DATA_OUT_1_6[21]\, DATA_OUT_1_6(20) => 
        \DATA_OUT_1_6[20]\, DATA_OUT_1_6(19) => 
        \DATA_OUT_1_6[19]\, DATA_OUT_1_6(18) => 
        \DATA_OUT_1_6[18]\, DATA_OUT_1_6(17) => 
        \DATA_OUT_1_6[17]\, DATA_OUT_1_6(16) => 
        \DATA_OUT_1_6[16]\, DATA_OUT_1_6(15) => 
        \DATA_OUT_1_6[15]\, DATA_OUT_1_6(14) => 
        \DATA_OUT_1_6[14]\, DATA_OUT_1_6(13) => 
        \DATA_OUT_1_6[13]\, DATA_OUT_1_6(12) => 
        \DATA_OUT_1_6[12]\, DATA_OUT_1_6(11) => 
        \DATA_OUT_1_6[11]\, DATA_OUT_1_6(10) => 
        \DATA_OUT_1_6[10]\, DATA_OUT_1_6(9) => \DATA_OUT_1_6[9]\, 
        DATA_OUT_1_6(8) => \DATA_OUT_1_6[8]\, DATA_OUT_1_6(7) => 
        \DATA_OUT_1_6[7]\, DATA_OUT_1_6(6) => \DATA_OUT_1_6[6]\, 
        DATA_OUT_1_6(5) => \DATA_OUT_1_6[5]\, DATA_OUT_1_6(4) => 
        \DATA_OUT_1_6[4]\, DATA_OUT_1_6(3) => \DATA_OUT_1_6[3]\, 
        DATA_OUT_1_6(2) => \DATA_OUT_1_6[2]\, DATA_OUT_1_6(1) => 
        \DATA_OUT_1_6[1]\, DATA_OUT_1_6(0) => \DATA_OUT_1_6[0]\, 
        DATA_OUT_1_7(25) => \DATA_OUT_1_7[25]\, DATA_OUT_1_7(24)
         => \DATA_OUT_1_7[24]\, DATA_OUT_1_7(23) => 
        \DATA_OUT_1_7[23]\, DATA_OUT_1_7(22) => 
        \DATA_OUT_1_7[22]\, DATA_OUT_1_7(21) => 
        \DATA_OUT_1_7[21]\, DATA_OUT_1_7(20) => 
        \DATA_OUT_1_7[20]\, DATA_OUT_1_7(19) => 
        \DATA_OUT_1_7[19]\, DATA_OUT_1_7(18) => 
        \DATA_OUT_1_7[18]\, DATA_OUT_1_7(17) => 
        \DATA_OUT_1_7[17]\, DATA_OUT_1_7(16) => 
        \DATA_OUT_1_7[16]\, DATA_OUT_1_7(15) => 
        \DATA_OUT_1_7[15]\, DATA_OUT_1_7(14) => 
        \DATA_OUT_1_7[14]\, DATA_OUT_1_7(13) => 
        \DATA_OUT_1_7[13]\, DATA_OUT_1_7(12) => 
        \DATA_OUT_1_7[12]\, DATA_OUT_1_7(11) => 
        \DATA_OUT_1_7[11]\, DATA_OUT_1_7(10) => 
        \DATA_OUT_1_7[10]\, DATA_OUT_1_7(9) => \DATA_OUT_1_7[9]\, 
        DATA_OUT_1_7(8) => \DATA_OUT_1_7[8]\, DATA_OUT_1_7(7) => 
        \DATA_OUT_1_7[7]\, DATA_OUT_1_7(6) => \DATA_OUT_1_7[6]\, 
        DATA_OUT_1_7(5) => \DATA_OUT_1_7[5]\, DATA_OUT_1_7(4) => 
        \DATA_OUT_1_7[4]\, DATA_OUT_1_7(3) => \DATA_OUT_1_7[3]\, 
        DATA_OUT_1_7(2) => \DATA_OUT_1_7[2]\, DATA_OUT_1_7(1) => 
        \DATA_OUT_1_7[1]\, DATA_OUT_1_7(0) => \DATA_OUT_1_7[0]\, 
        DATA_OUT_1_8(25) => \DATA_OUT_1_8[25]\, DATA_OUT_1_8(24)
         => \DATA_OUT_1_8[24]\, DATA_OUT_1_8(23) => 
        \DATA_OUT_1_8[23]\, DATA_OUT_1_8(22) => 
        \DATA_OUT_1_8[22]\, DATA_OUT_1_8(21) => 
        \DATA_OUT_1_8[21]\, DATA_OUT_1_8(20) => 
        \DATA_OUT_1_8[20]\, DATA_OUT_1_8(19) => 
        \DATA_OUT_1_8[19]\, DATA_OUT_1_8(18) => 
        \DATA_OUT_1_8[18]\, DATA_OUT_1_8(17) => 
        \DATA_OUT_1_8[17]\, DATA_OUT_1_8(16) => 
        \DATA_OUT_1_8[16]\, DATA_OUT_1_8(15) => 
        \DATA_OUT_1_8[15]\, DATA_OUT_1_8(14) => 
        \DATA_OUT_1_8[14]\, DATA_OUT_1_8(13) => 
        \DATA_OUT_1_8[13]\, DATA_OUT_1_8(12) => 
        \DATA_OUT_1_8[12]\, DATA_OUT_1_8(11) => 
        \DATA_OUT_1_8[11]\, DATA_OUT_1_8(10) => 
        \DATA_OUT_1_8[10]\, DATA_OUT_1_8(9) => \DATA_OUT_1_8[9]\, 
        DATA_OUT_1_8(8) => \DATA_OUT_1_8[8]\, DATA_OUT_1_8(7) => 
        \DATA_OUT_1_8[7]\, DATA_OUT_1_8(6) => \DATA_OUT_1_8[6]\, 
        DATA_OUT_1_8(5) => \DATA_OUT_1_8[5]\, DATA_OUT_1_8(4) => 
        \DATA_OUT_1_8[4]\, DATA_OUT_1_8(3) => \DATA_OUT_1_8[3]\, 
        DATA_OUT_1_8(2) => \DATA_OUT_1_8[2]\, DATA_OUT_1_8(1) => 
        \DATA_OUT_1_8[1]\, DATA_OUT_1_8(0) => \DATA_OUT_1_8[0]\, 
        DATA_OUT_1_9(25) => \DATA_OUT_1_9[25]\, DATA_OUT_1_9(24)
         => \DATA_OUT_1_9[24]\, DATA_OUT_1_9(23) => 
        \DATA_OUT_1_9[23]\, DATA_OUT_1_9(22) => 
        \DATA_OUT_1_9[22]\, DATA_OUT_1_9(21) => 
        \DATA_OUT_1_9[21]\, DATA_OUT_1_9(20) => 
        \DATA_OUT_1_9[20]\, DATA_OUT_1_9(19) => 
        \DATA_OUT_1_9[19]\, DATA_OUT_1_9(18) => 
        \DATA_OUT_1_9[18]\, DATA_OUT_1_9(17) => 
        \DATA_OUT_1_9[17]\, DATA_OUT_1_9(16) => 
        \DATA_OUT_1_9[16]\, DATA_OUT_1_9(15) => 
        \DATA_OUT_1_9[15]\, DATA_OUT_1_9(14) => 
        \DATA_OUT_1_9[14]\, DATA_OUT_1_9(13) => 
        \DATA_OUT_1_9[13]\, DATA_OUT_1_9(12) => 
        \DATA_OUT_1_9[12]\, DATA_OUT_1_9(11) => 
        \DATA_OUT_1_9[11]\, DATA_OUT_1_9(10) => 
        \DATA_OUT_1_9[10]\, DATA_OUT_1_9(9) => \DATA_OUT_1_9[9]\, 
        DATA_OUT_1_9(8) => \DATA_OUT_1_9[8]\, DATA_OUT_1_9(7) => 
        \DATA_OUT_1_9[7]\, DATA_OUT_1_9(6) => \DATA_OUT_1_9[6]\, 
        DATA_OUT_1_9(5) => \DATA_OUT_1_9[5]\, DATA_OUT_1_9(4) => 
        \DATA_OUT_1_9[4]\, DATA_OUT_1_9(3) => \DATA_OUT_1_9[3]\, 
        DATA_OUT_1_9(2) => \DATA_OUT_1_9[2]\, DATA_OUT_1_9(1) => 
        \DATA_OUT_1_9[1]\, DATA_OUT_1_9(0) => \DATA_OUT_1_9[0]\, 
        DATA_OUT_1_10(25) => \DATA_OUT_1_10[25]\, 
        DATA_OUT_1_10(24) => \DATA_OUT_1_10[24]\, 
        DATA_OUT_1_10(23) => \DATA_OUT_1_10[23]\, 
        DATA_OUT_1_10(22) => \DATA_OUT_1_10[22]\, 
        DATA_OUT_1_10(21) => \DATA_OUT_1_10[21]\, 
        DATA_OUT_1_10(20) => \DATA_OUT_1_10[20]\, 
        DATA_OUT_1_10(19) => \DATA_OUT_1_10[19]\, 
        DATA_OUT_1_10(18) => \DATA_OUT_1_10[18]\, 
        DATA_OUT_1_10(17) => \DATA_OUT_1_10[17]\, 
        DATA_OUT_1_10(16) => \DATA_OUT_1_10[16]\, 
        DATA_OUT_1_10(15) => \DATA_OUT_1_10[15]\, 
        DATA_OUT_1_10(14) => \DATA_OUT_1_10[14]\, 
        DATA_OUT_1_10(13) => \DATA_OUT_1_10[13]\, 
        DATA_OUT_1_10(12) => \DATA_OUT_1_10[12]\, 
        DATA_OUT_1_10(11) => \DATA_OUT_1_10[11]\, 
        DATA_OUT_1_10(10) => \DATA_OUT_1_10[10]\, 
        DATA_OUT_1_10(9) => \DATA_OUT_1_10[9]\, DATA_OUT_1_10(8)
         => \DATA_OUT_1_10[8]\, DATA_OUT_1_10(7) => 
        \DATA_OUT_1_10[7]\, DATA_OUT_1_10(6) => 
        \DATA_OUT_1_10[6]\, DATA_OUT_1_10(5) => 
        \DATA_OUT_1_10[5]\, DATA_OUT_1_10(4) => 
        \DATA_OUT_1_10[4]\, DATA_OUT_1_10(3) => 
        \DATA_OUT_1_10[3]\, DATA_OUT_1_10(2) => 
        \DATA_OUT_1_10[2]\, DATA_OUT_1_10(1) => 
        \DATA_OUT_1_10[1]\, DATA_OUT_1_10(0) => 
        \DATA_OUT_1_10[0]\, DATA_OUT_1_11(25) => 
        \DATA_OUT_1_11[25]\, DATA_OUT_1_11(24) => 
        \DATA_OUT_1_11[24]\, DATA_OUT_1_11(23) => 
        \DATA_OUT_1_11[23]\, DATA_OUT_1_11(22) => 
        \DATA_OUT_1_11[22]\, DATA_OUT_1_11(21) => 
        \DATA_OUT_1_11[21]\, DATA_OUT_1_11(20) => 
        \DATA_OUT_1_11[20]\, DATA_OUT_1_11(19) => 
        \DATA_OUT_1_11[19]\, DATA_OUT_1_11(18) => 
        \DATA_OUT_1_11[18]\, DATA_OUT_1_11(17) => 
        \DATA_OUT_1_11[17]\, DATA_OUT_1_11(16) => 
        \DATA_OUT_1_11[16]\, DATA_OUT_1_11(15) => 
        \DATA_OUT_1_11[15]\, DATA_OUT_1_11(14) => 
        \DATA_OUT_1_11[14]\, DATA_OUT_1_11(13) => 
        \DATA_OUT_1_11[13]\, DATA_OUT_1_11(12) => 
        \DATA_OUT_1_11[12]\, DATA_OUT_1_11(11) => 
        \DATA_OUT_1_11[11]\, DATA_OUT_1_11(10) => 
        \DATA_OUT_1_11[10]\, DATA_OUT_1_11(9) => 
        \DATA_OUT_1_11[9]\, DATA_OUT_1_11(8) => 
        \DATA_OUT_1_11[8]\, DATA_OUT_1_11(7) => 
        \DATA_OUT_1_11[7]\, DATA_OUT_1_11(6) => 
        \DATA_OUT_1_11[6]\, DATA_OUT_1_11(5) => 
        \DATA_OUT_1_11[5]\, DATA_OUT_1_11(4) => 
        \DATA_OUT_1_11[4]\, DATA_OUT_1_11(3) => 
        \DATA_OUT_1_11[3]\, DATA_OUT_1_11(2) => 
        \DATA_OUT_1_11[2]\, DATA_OUT_1_11(1) => 
        \DATA_OUT_1_11[1]\, DATA_OUT_1_11(0) => 
        \DATA_OUT_1_11[0]\, DATA_OUT_1_12(25) => 
        \DATA_OUT_1_12[25]\, DATA_OUT_1_12(24) => 
        \DATA_OUT_1_12[24]\, DATA_OUT_1_12(23) => 
        \DATA_OUT_1_12[23]\, DATA_OUT_1_12(22) => 
        \DATA_OUT_1_12[22]\, DATA_OUT_1_12(21) => 
        \DATA_OUT_1_12[21]\, DATA_OUT_1_12(20) => 
        \DATA_OUT_1_12[20]\, DATA_OUT_1_12(19) => 
        \DATA_OUT_1_12[19]\, DATA_OUT_1_12(18) => 
        \DATA_OUT_1_12[18]\, DATA_OUT_1_12(17) => 
        \DATA_OUT_1_12[17]\, DATA_OUT_1_12(16) => 
        \DATA_OUT_1_12[16]\, DATA_OUT_1_12(15) => 
        \DATA_OUT_1_12[15]\, DATA_OUT_1_12(14) => 
        \DATA_OUT_1_12[14]\, DATA_OUT_1_12(13) => 
        \DATA_OUT_1_12[13]\, DATA_OUT_1_12(12) => 
        \DATA_OUT_1_12[12]\, DATA_OUT_1_12(11) => 
        \DATA_OUT_1_12[11]\, DATA_OUT_1_12(10) => 
        \DATA_OUT_1_12[10]\, DATA_OUT_1_12(9) => 
        \DATA_OUT_1_12[9]\, DATA_OUT_1_12(8) => 
        \DATA_OUT_1_12[8]\, DATA_OUT_1_12(7) => 
        \DATA_OUT_1_12[7]\, DATA_OUT_1_12(6) => 
        \DATA_OUT_1_12[6]\, DATA_OUT_1_12(5) => 
        \DATA_OUT_1_12[5]\, DATA_OUT_1_12(4) => 
        \DATA_OUT_1_12[4]\, DATA_OUT_1_12(3) => 
        \DATA_OUT_1_12[3]\, DATA_OUT_1_12(2) => 
        \DATA_OUT_1_12[2]\, DATA_OUT_1_12(1) => 
        \DATA_OUT_1_12[1]\, DATA_OUT_1_12(0) => 
        \DATA_OUT_1_12[0]\, DATA_OUT_1_13(25) => 
        \DATA_OUT_1_13[25]\, DATA_OUT_1_13(24) => 
        \DATA_OUT_1_13[24]\, DATA_OUT_1_13(23) => 
        \DATA_OUT_1_13[23]\, DATA_OUT_1_13(22) => 
        \DATA_OUT_1_13[22]\, DATA_OUT_1_13(21) => 
        \DATA_OUT_1_13[21]\, DATA_OUT_1_13(20) => 
        \DATA_OUT_1_13[20]\, DATA_OUT_1_13(19) => 
        \DATA_OUT_1_13[19]\, DATA_OUT_1_13(18) => 
        \DATA_OUT_1_13[18]\, DATA_OUT_1_13(17) => 
        \DATA_OUT_1_13[17]\, DATA_OUT_1_13(16) => 
        \DATA_OUT_1_13[16]\, DATA_OUT_1_13(15) => 
        \DATA_OUT_1_13[15]\, DATA_OUT_1_13(14) => 
        \DATA_OUT_1_13[14]\, DATA_OUT_1_13(13) => 
        \DATA_OUT_1_13[13]\, DATA_OUT_1_13(12) => 
        \DATA_OUT_1_13[12]\, DATA_OUT_1_13(11) => 
        \DATA_OUT_1_13[11]\, DATA_OUT_1_13(10) => 
        \DATA_OUT_1_13[10]\, DATA_OUT_1_13(9) => 
        \DATA_OUT_1_13[9]\, DATA_OUT_1_13(8) => 
        \DATA_OUT_1_13[8]\, DATA_OUT_1_13(7) => 
        \DATA_OUT_1_13[7]\, DATA_OUT_1_13(6) => 
        \DATA_OUT_1_13[6]\, DATA_OUT_1_13(5) => 
        \DATA_OUT_1_13[5]\, DATA_OUT_1_13(4) => 
        \DATA_OUT_1_13[4]\, DATA_OUT_1_13(3) => 
        \DATA_OUT_1_13[3]\, DATA_OUT_1_13(2) => 
        \DATA_OUT_1_13[2]\, DATA_OUT_1_13(1) => 
        \DATA_OUT_1_13[1]\, DATA_OUT_1_13(0) => 
        \DATA_OUT_1_13[0]\, DATA_OUT_1_14(25) => 
        \DATA_OUT_1_14[25]\, DATA_OUT_1_14(24) => 
        \DATA_OUT_1_14[24]\, DATA_OUT_1_14(23) => 
        \DATA_OUT_1_14[23]\, DATA_OUT_1_14(22) => 
        \DATA_OUT_1_14[22]\, DATA_OUT_1_14(21) => 
        \DATA_OUT_1_14[21]\, DATA_OUT_1_14(20) => 
        \DATA_OUT_1_14[20]\, DATA_OUT_1_14(19) => 
        \DATA_OUT_1_14[19]\, DATA_OUT_1_14(18) => 
        \DATA_OUT_1_14[18]\, DATA_OUT_1_14(17) => 
        \DATA_OUT_1_14[17]\, DATA_OUT_1_14(16) => 
        \DATA_OUT_1_14[16]\, DATA_OUT_1_14(15) => 
        \DATA_OUT_1_14[15]\, DATA_OUT_1_14(14) => 
        \DATA_OUT_1_14[14]\, DATA_OUT_1_14(13) => 
        \DATA_OUT_1_14[13]\, DATA_OUT_1_14(12) => 
        \DATA_OUT_1_14[12]\, DATA_OUT_1_14(11) => 
        \DATA_OUT_1_14[11]\, DATA_OUT_1_14(10) => 
        \DATA_OUT_1_14[10]\, DATA_OUT_1_14(9) => 
        \DATA_OUT_1_14[9]\, DATA_OUT_1_14(8) => 
        \DATA_OUT_1_14[8]\, DATA_OUT_1_14(7) => 
        \DATA_OUT_1_14[7]\, DATA_OUT_1_14(6) => 
        \DATA_OUT_1_14[6]\, DATA_OUT_1_14(5) => 
        \DATA_OUT_1_14[5]\, DATA_OUT_1_14(4) => 
        \DATA_OUT_1_14[4]\, DATA_OUT_1_14(3) => 
        \DATA_OUT_1_14[3]\, DATA_OUT_1_14(2) => 
        \DATA_OUT_1_14[2]\, DATA_OUT_1_14(1) => 
        \DATA_OUT_1_14[1]\, DATA_OUT_1_14(0) => 
        \DATA_OUT_1_14[0]\, DATA_OUT_1_15(25) => 
        \DATA_OUT_1_15[25]\, DATA_OUT_1_15(24) => 
        \DATA_OUT_1_15[24]\, DATA_OUT_1_15(23) => 
        \DATA_OUT_1_15[23]\, DATA_OUT_1_15(22) => 
        \DATA_OUT_1_15[22]\, DATA_OUT_1_15(21) => 
        \DATA_OUT_1_15[21]\, DATA_OUT_1_15(20) => 
        \DATA_OUT_1_15[20]\, DATA_OUT_1_15(19) => 
        \DATA_OUT_1_15[19]\, DATA_OUT_1_15(18) => 
        \DATA_OUT_1_15[18]\, DATA_OUT_1_15(17) => 
        \DATA_OUT_1_15[17]\, DATA_OUT_1_15(16) => 
        \DATA_OUT_1_15[16]\, DATA_OUT_1_15(15) => 
        \DATA_OUT_1_15[15]\, DATA_OUT_1_15(14) => 
        \DATA_OUT_1_15[14]\, DATA_OUT_1_15(13) => 
        \DATA_OUT_1_15[13]\, DATA_OUT_1_15(12) => 
        \DATA_OUT_1_15[12]\, DATA_OUT_1_15(11) => 
        \DATA_OUT_1_15[11]\, DATA_OUT_1_15(10) => 
        \DATA_OUT_1_15[10]\, DATA_OUT_1_15(9) => 
        \DATA_OUT_1_15[9]\, DATA_OUT_1_15(8) => 
        \DATA_OUT_1_15[8]\, DATA_OUT_1_15(7) => 
        \DATA_OUT_1_15[7]\, DATA_OUT_1_15(6) => 
        \DATA_OUT_1_15[6]\, DATA_OUT_1_15(5) => 
        \DATA_OUT_1_15[5]\, DATA_OUT_1_15(4) => 
        \DATA_OUT_1_15[4]\, DATA_OUT_1_15(3) => 
        \DATA_OUT_1_15[3]\, DATA_OUT_1_15(2) => 
        \DATA_OUT_1_15[2]\, DATA_OUT_1_15(1) => 
        \DATA_OUT_1_15[1]\, DATA_OUT_1_15(0) => 
        \DATA_OUT_1_15[0]\, DATA_OUT_1_16(25) => 
        \DATA_OUT_1_16[25]\, DATA_OUT_1_16(24) => 
        \DATA_OUT_1_16[24]\, DATA_OUT_1_16(23) => 
        \DATA_OUT_1_16[23]\, DATA_OUT_1_16(22) => 
        \DATA_OUT_1_16[22]\, DATA_OUT_1_16(21) => 
        \DATA_OUT_1_16[21]\, DATA_OUT_1_16(20) => 
        \DATA_OUT_1_16[20]\, DATA_OUT_1_16(19) => 
        \DATA_OUT_1_16[19]\, DATA_OUT_1_16(18) => 
        \DATA_OUT_1_16[18]\, DATA_OUT_1_16(17) => 
        \DATA_OUT_1_16[17]\, DATA_OUT_1_16(16) => 
        \DATA_OUT_1_16[16]\, DATA_OUT_1_16(15) => 
        \DATA_OUT_1_16[15]\, DATA_OUT_1_16(14) => 
        \DATA_OUT_1_16[14]\, DATA_OUT_1_16(13) => 
        \DATA_OUT_1_16[13]\, DATA_OUT_1_16(12) => 
        \DATA_OUT_1_16[12]\, DATA_OUT_1_16(11) => 
        \DATA_OUT_1_16[11]\, DATA_OUT_1_16(10) => 
        \DATA_OUT_1_16[10]\, DATA_OUT_1_16(9) => 
        \DATA_OUT_1_16[9]\, DATA_OUT_1_16(8) => 
        \DATA_OUT_1_16[8]\, DATA_OUT_1_16(7) => 
        \DATA_OUT_1_16[7]\, DATA_OUT_1_16(6) => 
        \DATA_OUT_1_16[6]\, DATA_OUT_1_16(5) => 
        \DATA_OUT_1_16[5]\, DATA_OUT_1_16(4) => 
        \DATA_OUT_1_16[4]\, DATA_OUT_1_16(3) => 
        \DATA_OUT_1_16[3]\, DATA_OUT_1_16(2) => 
        \DATA_OUT_1_16[2]\, DATA_OUT_1_16(1) => 
        \DATA_OUT_1_16[1]\, DATA_OUT_1_16(0) => 
        \DATA_OUT_1_16[0]\, DATA_OUT_1_17(25) => 
        \DATA_OUT_1_17[25]\, DATA_OUT_1_17(24) => 
        \DATA_OUT_1_17[24]\, DATA_OUT_1_17(23) => 
        \DATA_OUT_1_17[23]\, DATA_OUT_1_17(22) => 
        \DATA_OUT_1_17[22]\, DATA_OUT_1_17(21) => 
        \DATA_OUT_1_17[21]\, DATA_OUT_1_17(20) => 
        \DATA_OUT_1_17[20]\, DATA_OUT_1_17(19) => 
        \DATA_OUT_1_17[19]\, DATA_OUT_1_17(18) => 
        \DATA_OUT_1_17[18]\, DATA_OUT_1_17(17) => 
        \DATA_OUT_1_17[17]\, DATA_OUT_1_17(16) => 
        \DATA_OUT_1_17[16]\, DATA_OUT_1_17(15) => 
        \DATA_OUT_1_17[15]\, DATA_OUT_1_17(14) => 
        \DATA_OUT_1_17[14]\, DATA_OUT_1_17(13) => 
        \DATA_OUT_1_17[13]\, DATA_OUT_1_17(12) => 
        \DATA_OUT_1_17[12]\, DATA_OUT_1_17(11) => 
        \DATA_OUT_1_17[11]\, DATA_OUT_1_17(10) => 
        \DATA_OUT_1_17[10]\, DATA_OUT_1_17(9) => 
        \DATA_OUT_1_17[9]\, DATA_OUT_1_17(8) => 
        \DATA_OUT_1_17[8]\, DATA_OUT_1_17(7) => 
        \DATA_OUT_1_17[7]\, DATA_OUT_1_17(6) => 
        \DATA_OUT_1_17[6]\, DATA_OUT_1_17(5) => 
        \DATA_OUT_1_17[5]\, DATA_OUT_1_17(4) => 
        \DATA_OUT_1_17[4]\, DATA_OUT_1_17(3) => 
        \DATA_OUT_1_17[3]\, DATA_OUT_1_17(2) => 
        \DATA_OUT_1_17[2]\, DATA_OUT_1_17(1) => 
        \DATA_OUT_1_17[1]\, DATA_OUT_1_17(0) => 
        \DATA_OUT_1_17[0]\, DATA_OUT_1_18(25) => 
        \DATA_OUT_1_18[25]\, DATA_OUT_1_18(24) => 
        \DATA_OUT_1_18[24]\, DATA_OUT_1_18(23) => 
        \DATA_OUT_1_18[23]\, DATA_OUT_1_18(22) => 
        \DATA_OUT_1_18[22]\, DATA_OUT_1_18(21) => 
        \DATA_OUT_1_18[21]\, DATA_OUT_1_18(20) => 
        \DATA_OUT_1_18[20]\, DATA_OUT_1_18(19) => 
        \DATA_OUT_1_18[19]\, DATA_OUT_1_18(18) => 
        \DATA_OUT_1_18[18]\, DATA_OUT_1_18(17) => 
        \DATA_OUT_1_18[17]\, DATA_OUT_1_18(16) => 
        \DATA_OUT_1_18[16]\, DATA_OUT_1_18(15) => 
        \DATA_OUT_1_18[15]\, DATA_OUT_1_18(14) => 
        \DATA_OUT_1_18[14]\, DATA_OUT_1_18(13) => 
        \DATA_OUT_1_18[13]\, DATA_OUT_1_18(12) => 
        \DATA_OUT_1_18[12]\, DATA_OUT_1_18(11) => 
        \DATA_OUT_1_18[11]\, DATA_OUT_1_18(10) => 
        \DATA_OUT_1_18[10]\, DATA_OUT_1_18(9) => 
        \DATA_OUT_1_18[9]\, DATA_OUT_1_18(8) => 
        \DATA_OUT_1_18[8]\, DATA_OUT_1_18(7) => 
        \DATA_OUT_1_18[7]\, DATA_OUT_1_18(6) => 
        \DATA_OUT_1_18[6]\, DATA_OUT_1_18(5) => 
        \DATA_OUT_1_18[5]\, DATA_OUT_1_18(4) => 
        \DATA_OUT_1_18[4]\, DATA_OUT_1_18(3) => 
        \DATA_OUT_1_18[3]\, DATA_OUT_1_18(2) => 
        \DATA_OUT_1_18[2]\, DATA_OUT_1_18(1) => 
        \DATA_OUT_1_18[1]\, DATA_OUT_1_18(0) => 
        \DATA_OUT_1_18[0]\, DATA_OUT_1_19(25) => 
        \DATA_OUT_1_19[25]\, DATA_OUT_1_19(24) => 
        \DATA_OUT_1_19[24]\, DATA_OUT_1_19(23) => 
        \DATA_OUT_1_19[23]\, DATA_OUT_1_19(22) => 
        \DATA_OUT_1_19[22]\, DATA_OUT_1_19(21) => 
        \DATA_OUT_1_19[21]\, DATA_OUT_1_19(20) => 
        \DATA_OUT_1_19[20]\, DATA_OUT_1_19(19) => 
        \DATA_OUT_1_19[19]\, DATA_OUT_1_19(18) => 
        \DATA_OUT_1_19[18]\, DATA_OUT_1_19(17) => 
        \DATA_OUT_1_19[17]\, DATA_OUT_1_19(16) => 
        \DATA_OUT_1_19[16]\, DATA_OUT_1_19(15) => 
        \DATA_OUT_1_19[15]\, DATA_OUT_1_19(14) => 
        \DATA_OUT_1_19[14]\, DATA_OUT_1_19(13) => 
        \DATA_OUT_1_19[13]\, DATA_OUT_1_19(12) => 
        \DATA_OUT_1_19[12]\, DATA_OUT_1_19(11) => 
        \DATA_OUT_1_19[11]\, DATA_OUT_1_19(10) => 
        \DATA_OUT_1_19[10]\, DATA_OUT_1_19(9) => 
        \DATA_OUT_1_19[9]\, DATA_OUT_1_19(8) => 
        \DATA_OUT_1_19[8]\, DATA_OUT_1_19(7) => 
        \DATA_OUT_1_19[7]\, DATA_OUT_1_19(6) => 
        \DATA_OUT_1_19[6]\, DATA_OUT_1_19(5) => 
        \DATA_OUT_1_19[5]\, DATA_OUT_1_19(4) => 
        \DATA_OUT_1_19[4]\, DATA_OUT_1_19(3) => 
        \DATA_OUT_1_19[3]\, DATA_OUT_1_19(2) => 
        \DATA_OUT_1_19[2]\, DATA_OUT_1_19(1) => 
        \DATA_OUT_1_19[1]\, DATA_OUT_1_19(0) => 
        \DATA_OUT_1_19[0]\, DATA_OUT_1_20(25) => 
        \DATA_OUT_1_20[25]\, DATA_OUT_1_20(24) => 
        \DATA_OUT_1_20[24]\, DATA_OUT_1_20(23) => 
        \DATA_OUT_1_20[23]\, DATA_OUT_1_20(22) => 
        \DATA_OUT_1_20[22]\, DATA_OUT_1_20(21) => 
        \DATA_OUT_1_20[21]\, DATA_OUT_1_20(20) => 
        \DATA_OUT_1_20[20]\, DATA_OUT_1_20(19) => 
        \DATA_OUT_1_20[19]\, DATA_OUT_1_20(18) => 
        \DATA_OUT_1_20[18]\, DATA_OUT_1_20(17) => 
        \DATA_OUT_1_20[17]\, DATA_OUT_1_20(16) => 
        \DATA_OUT_1_20[16]\, DATA_OUT_1_20(15) => 
        \DATA_OUT_1_20[15]\, DATA_OUT_1_20(14) => 
        \DATA_OUT_1_20[14]\, DATA_OUT_1_20(13) => 
        \DATA_OUT_1_20[13]\, DATA_OUT_1_20(12) => 
        \DATA_OUT_1_20[12]\, DATA_OUT_1_20(11) => 
        \DATA_OUT_1_20[11]\, DATA_OUT_1_20(10) => 
        \DATA_OUT_1_20[10]\, DATA_OUT_1_20(9) => 
        \DATA_OUT_1_20[9]\, DATA_OUT_1_20(8) => 
        \DATA_OUT_1_20[8]\, DATA_OUT_1_20(7) => 
        \DATA_OUT_1_20[7]\, DATA_OUT_1_20(6) => 
        \DATA_OUT_1_20[6]\, DATA_OUT_1_20(5) => 
        \DATA_OUT_1_20[5]\, DATA_OUT_1_20(4) => 
        \DATA_OUT_1_20[4]\, DATA_OUT_1_20(3) => 
        \DATA_OUT_1_20[3]\, DATA_OUT_1_20(2) => 
        \DATA_OUT_1_20[2]\, DATA_OUT_1_20(1) => 
        \DATA_OUT_1_20[1]\, DATA_OUT_1_20(0) => 
        \DATA_OUT_1_20[0]\, DATA_OUT_1_21(25) => 
        \DATA_OUT_1_21[25]\, DATA_OUT_1_21(24) => 
        \DATA_OUT_1_21[24]\, DATA_OUT_1_21(23) => 
        \DATA_OUT_1_21[23]\, DATA_OUT_1_21(22) => 
        \DATA_OUT_1_21[22]\, DATA_OUT_1_21(21) => 
        \DATA_OUT_1_21[21]\, DATA_OUT_1_21(20) => 
        \DATA_OUT_1_21[20]\, DATA_OUT_1_21(19) => 
        \DATA_OUT_1_21[19]\, DATA_OUT_1_21(18) => 
        \DATA_OUT_1_21[18]\, DATA_OUT_1_21(17) => 
        \DATA_OUT_1_21[17]\, DATA_OUT_1_21(16) => 
        \DATA_OUT_1_21[16]\, DATA_OUT_1_21(15) => 
        \DATA_OUT_1_21[15]\, DATA_OUT_1_21(14) => 
        \DATA_OUT_1_21[14]\, DATA_OUT_1_21(13) => 
        \DATA_OUT_1_21[13]\, DATA_OUT_1_21(12) => 
        \DATA_OUT_1_21[12]\, DATA_OUT_1_21(11) => 
        \DATA_OUT_1_21[11]\, DATA_OUT_1_21(10) => 
        \DATA_OUT_1_21[10]\, DATA_OUT_1_21(9) => 
        \DATA_OUT_1_21[9]\, DATA_OUT_1_21(8) => 
        \DATA_OUT_1_21[8]\, DATA_OUT_1_21(7) => 
        \DATA_OUT_1_21[7]\, DATA_OUT_1_21(6) => 
        \DATA_OUT_1_21[6]\, DATA_OUT_1_21(5) => 
        \DATA_OUT_1_21[5]\, DATA_OUT_1_21(4) => 
        \DATA_OUT_1_21[4]\, DATA_OUT_1_21(3) => 
        \DATA_OUT_1_21[3]\, DATA_OUT_1_21(2) => 
        \DATA_OUT_1_21[2]\, DATA_OUT_1_21(1) => 
        \DATA_OUT_1_21[1]\, DATA_OUT_1_21(0) => 
        \DATA_OUT_1_21[0]\, DATA_OUT_1_22(25) => 
        \DATA_OUT_1_22[25]\, DATA_OUT_1_22(24) => 
        \DATA_OUT_1_22[24]\, DATA_OUT_1_22(23) => 
        \DATA_OUT_1_22[23]\, DATA_OUT_1_22(22) => 
        \DATA_OUT_1_22[22]\, DATA_OUT_1_22(21) => 
        \DATA_OUT_1_22[21]\, DATA_OUT_1_22(20) => 
        \DATA_OUT_1_22[20]\, DATA_OUT_1_22(19) => 
        \DATA_OUT_1_22[19]\, DATA_OUT_1_22(18) => 
        \DATA_OUT_1_22[18]\, DATA_OUT_1_22(17) => 
        \DATA_OUT_1_22[17]\, DATA_OUT_1_22(16) => 
        \DATA_OUT_1_22[16]\, DATA_OUT_1_22(15) => 
        \DATA_OUT_1_22[15]\, DATA_OUT_1_22(14) => 
        \DATA_OUT_1_22[14]\, DATA_OUT_1_22(13) => 
        \DATA_OUT_1_22[13]\, DATA_OUT_1_22(12) => 
        \DATA_OUT_1_22[12]\, DATA_OUT_1_22(11) => 
        \DATA_OUT_1_22[11]\, DATA_OUT_1_22(10) => 
        \DATA_OUT_1_22[10]\, DATA_OUT_1_22(9) => 
        \DATA_OUT_1_22[9]\, DATA_OUT_1_22(8) => 
        \DATA_OUT_1_22[8]\, DATA_OUT_1_22(7) => 
        \DATA_OUT_1_22[7]\, DATA_OUT_1_22(6) => 
        \DATA_OUT_1_22[6]\, DATA_OUT_1_22(5) => 
        \DATA_OUT_1_22[5]\, DATA_OUT_1_22(4) => 
        \DATA_OUT_1_22[4]\, DATA_OUT_1_22(3) => 
        \DATA_OUT_1_22[3]\, DATA_OUT_1_22(2) => 
        \DATA_OUT_1_22[2]\, DATA_OUT_1_22(1) => 
        \DATA_OUT_1_22[1]\, DATA_OUT_1_22(0) => 
        \DATA_OUT_1_22[0]\, DATA_OUT_1_23(25) => 
        \DATA_OUT_1_23[25]\, DATA_OUT_1_23(24) => 
        \DATA_OUT_1_23[24]\, DATA_OUT_1_23(23) => 
        \DATA_OUT_1_23[23]\, DATA_OUT_1_23(22) => 
        \DATA_OUT_1_23[22]\, DATA_OUT_1_23(21) => 
        \DATA_OUT_1_23[21]\, DATA_OUT_1_23(20) => 
        \DATA_OUT_1_23[20]\, DATA_OUT_1_23(19) => 
        \DATA_OUT_1_23[19]\, DATA_OUT_1_23(18) => 
        \DATA_OUT_1_23[18]\, DATA_OUT_1_23(17) => 
        \DATA_OUT_1_23[17]\, DATA_OUT_1_23(16) => 
        \DATA_OUT_1_23[16]\, DATA_OUT_1_23(15) => 
        \DATA_OUT_1_23[15]\, DATA_OUT_1_23(14) => 
        \DATA_OUT_1_23[14]\, DATA_OUT_1_23(13) => 
        \DATA_OUT_1_23[13]\, DATA_OUT_1_23(12) => 
        \DATA_OUT_1_23[12]\, DATA_OUT_1_23(11) => 
        \DATA_OUT_1_23[11]\, DATA_OUT_1_23(10) => 
        \DATA_OUT_1_23[10]\, DATA_OUT_1_23(9) => 
        \DATA_OUT_1_23[9]\, DATA_OUT_1_23(8) => 
        \DATA_OUT_1_23[8]\, DATA_OUT_1_23(7) => 
        \DATA_OUT_1_23[7]\, DATA_OUT_1_23(6) => 
        \DATA_OUT_1_23[6]\, DATA_OUT_1_23(5) => 
        \DATA_OUT_1_23[5]\, DATA_OUT_1_23(4) => 
        \DATA_OUT_1_23[4]\, DATA_OUT_1_23(3) => 
        \DATA_OUT_1_23[3]\, DATA_OUT_1_23(2) => 
        \DATA_OUT_1_23[2]\, DATA_OUT_1_23(1) => 
        \DATA_OUT_1_23[1]\, DATA_OUT_1_23(0) => 
        \DATA_OUT_1_23[0]\, DATA_OUT_1_24(25) => 
        \DATA_OUT_1_24[25]\, DATA_OUT_1_24(24) => 
        \DATA_OUT_1_24[24]\, DATA_OUT_1_24(23) => 
        \DATA_OUT_1_24[23]\, DATA_OUT_1_24(22) => 
        \DATA_OUT_1_24[22]\, DATA_OUT_1_24(21) => 
        \DATA_OUT_1_24[21]\, DATA_OUT_1_24(20) => 
        \DATA_OUT_1_24[20]\, DATA_OUT_1_24(19) => 
        \DATA_OUT_1_24[19]\, DATA_OUT_1_24(18) => 
        \DATA_OUT_1_24[18]\, DATA_OUT_1_24(17) => 
        \DATA_OUT_1_24[17]\, DATA_OUT_1_24(16) => 
        \DATA_OUT_1_24[16]\, DATA_OUT_1_24(15) => 
        \DATA_OUT_1_24[15]\, DATA_OUT_1_24(14) => 
        \DATA_OUT_1_24[14]\, DATA_OUT_1_24(13) => 
        \DATA_OUT_1_24[13]\, DATA_OUT_1_24(12) => 
        \DATA_OUT_1_24[12]\, DATA_OUT_1_24(11) => 
        \DATA_OUT_1_24[11]\, DATA_OUT_1_24(10) => 
        \DATA_OUT_1_24[10]\, DATA_OUT_1_24(9) => 
        \DATA_OUT_1_24[9]\, DATA_OUT_1_24(8) => 
        \DATA_OUT_1_24[8]\, DATA_OUT_1_24(7) => 
        \DATA_OUT_1_24[7]\, DATA_OUT_1_24(6) => 
        \DATA_OUT_1_24[6]\, DATA_OUT_1_24(5) => 
        \DATA_OUT_1_24[5]\, DATA_OUT_1_24(4) => 
        \DATA_OUT_1_24[4]\, DATA_OUT_1_24(3) => 
        \DATA_OUT_1_24[3]\, DATA_OUT_1_24(2) => 
        \DATA_OUT_1_24[2]\, DATA_OUT_1_24(1) => 
        \DATA_OUT_1_24[1]\, DATA_OUT_1_24(0) => 
        \DATA_OUT_1_24[0]\, DATA_OUT_1_25(25) => 
        \DATA_OUT_1_25[25]\, DATA_OUT_1_25(24) => 
        \DATA_OUT_1_25[24]\, DATA_OUT_1_25(23) => 
        \DATA_OUT_1_25[23]\, DATA_OUT_1_25(22) => 
        \DATA_OUT_1_25[22]\, DATA_OUT_1_25(21) => 
        \DATA_OUT_1_25[21]\, DATA_OUT_1_25(20) => 
        \DATA_OUT_1_25[20]\, DATA_OUT_1_25(19) => 
        \DATA_OUT_1_25[19]\, DATA_OUT_1_25(18) => 
        \DATA_OUT_1_25[18]\, DATA_OUT_1_25(17) => 
        \DATA_OUT_1_25[17]\, DATA_OUT_1_25(16) => 
        \DATA_OUT_1_25[16]\, DATA_OUT_1_25(15) => 
        \DATA_OUT_1_25[15]\, DATA_OUT_1_25(14) => 
        \DATA_OUT_1_25[14]\, DATA_OUT_1_25(13) => 
        \DATA_OUT_1_25[13]\, DATA_OUT_1_25(12) => 
        \DATA_OUT_1_25[12]\, DATA_OUT_1_25(11) => 
        \DATA_OUT_1_25[11]\, DATA_OUT_1_25(10) => 
        \DATA_OUT_1_25[10]\, DATA_OUT_1_25(9) => 
        \DATA_OUT_1_25[9]\, DATA_OUT_1_25(8) => 
        \DATA_OUT_1_25[8]\, DATA_OUT_1_25(7) => 
        \DATA_OUT_1_25[7]\, DATA_OUT_1_25(6) => 
        \DATA_OUT_1_25[6]\, DATA_OUT_1_25(5) => 
        \DATA_OUT_1_25[5]\, DATA_OUT_1_25(4) => 
        \DATA_OUT_1_25[4]\, DATA_OUT_1_25(3) => 
        \DATA_OUT_1_25[3]\, DATA_OUT_1_25(2) => 
        \DATA_OUT_1_25[2]\, DATA_OUT_1_25(1) => 
        \DATA_OUT_1_25[1]\, DATA_OUT_1_25(0) => 
        \DATA_OUT_1_25[0]\, DATA_OUT_1_26(25) => 
        \DATA_OUT_1_26[25]\, DATA_OUT_1_26(24) => 
        \DATA_OUT_1_26[24]\, DATA_OUT_1_26(23) => 
        \DATA_OUT_1_26[23]\, DATA_OUT_1_26(22) => 
        \DATA_OUT_1_26[22]\, DATA_OUT_1_26(21) => 
        \DATA_OUT_1_26[21]\, DATA_OUT_1_26(20) => 
        \DATA_OUT_1_26[20]\, DATA_OUT_1_26(19) => 
        \DATA_OUT_1_26[19]\, DATA_OUT_1_26(18) => 
        \DATA_OUT_1_26[18]\, DATA_OUT_1_26(17) => 
        \DATA_OUT_1_26[17]\, DATA_OUT_1_26(16) => 
        \DATA_OUT_1_26[16]\, DATA_OUT_1_26(15) => 
        \DATA_OUT_1_26[15]\, DATA_OUT_1_26(14) => 
        \DATA_OUT_1_26[14]\, DATA_OUT_1_26(13) => 
        \DATA_OUT_1_26[13]\, DATA_OUT_1_26(12) => 
        \DATA_OUT_1_26[12]\, DATA_OUT_1_26(11) => 
        \DATA_OUT_1_26[11]\, DATA_OUT_1_26(10) => 
        \DATA_OUT_1_26[10]\, DATA_OUT_1_26(9) => 
        \DATA_OUT_1_26[9]\, DATA_OUT_1_26(8) => 
        \DATA_OUT_1_26[8]\, DATA_OUT_1_26(7) => 
        \DATA_OUT_1_26[7]\, DATA_OUT_1_26(6) => 
        \DATA_OUT_1_26[6]\, DATA_OUT_1_26(5) => 
        \DATA_OUT_1_26[5]\, DATA_OUT_1_26(4) => 
        \DATA_OUT_1_26[4]\, DATA_OUT_1_26(3) => 
        \DATA_OUT_1_26[3]\, DATA_OUT_1_26(2) => 
        \DATA_OUT_1_26[2]\, DATA_OUT_1_26(1) => 
        \DATA_OUT_1_26[1]\, DATA_OUT_1_26(0) => 
        \DATA_OUT_1_26[0]\, DATA_OUT_1_27(25) => 
        \DATA_OUT_1_27[25]\, DATA_OUT_1_27(24) => 
        \DATA_OUT_1_27[24]\, DATA_OUT_1_27(23) => 
        \DATA_OUT_1_27[23]\, DATA_OUT_1_27(22) => 
        \DATA_OUT_1_27[22]\, DATA_OUT_1_27(21) => 
        \DATA_OUT_1_27[21]\, DATA_OUT_1_27(20) => 
        \DATA_OUT_1_27[20]\, DATA_OUT_1_27(19) => 
        \DATA_OUT_1_27[19]\, DATA_OUT_1_27(18) => 
        \DATA_OUT_1_27[18]\, DATA_OUT_1_27(17) => 
        \DATA_OUT_1_27[17]\, DATA_OUT_1_27(16) => 
        \DATA_OUT_1_27[16]\, DATA_OUT_1_27(15) => 
        \DATA_OUT_1_27[15]\, DATA_OUT_1_27(14) => 
        \DATA_OUT_1_27[14]\, DATA_OUT_1_27(13) => 
        \DATA_OUT_1_27[13]\, DATA_OUT_1_27(12) => 
        \DATA_OUT_1_27[12]\, DATA_OUT_1_27(11) => 
        \DATA_OUT_1_27[11]\, DATA_OUT_1_27(10) => 
        \DATA_OUT_1_27[10]\, DATA_OUT_1_27(9) => 
        \DATA_OUT_1_27[9]\, DATA_OUT_1_27(8) => 
        \DATA_OUT_1_27[8]\, DATA_OUT_1_27(7) => 
        \DATA_OUT_1_27[7]\, DATA_OUT_1_27(6) => 
        \DATA_OUT_1_27[6]\, DATA_OUT_1_27(5) => 
        \DATA_OUT_1_27[5]\, DATA_OUT_1_27(4) => 
        \DATA_OUT_1_27[4]\, DATA_OUT_1_27(3) => 
        \DATA_OUT_1_27[3]\, DATA_OUT_1_27(2) => 
        \DATA_OUT_1_27[2]\, DATA_OUT_1_27(1) => 
        \DATA_OUT_1_27[1]\, DATA_OUT_1_27(0) => 
        \DATA_OUT_1_27[0]\, DATA_OUT_1_28(25) => 
        \DATA_OUT_1_28[25]\, DATA_OUT_1_28(24) => 
        \DATA_OUT_1_28[24]\, DATA_OUT_1_28(23) => 
        \DATA_OUT_1_28[23]\, DATA_OUT_1_28(22) => 
        \DATA_OUT_1_28[22]\, DATA_OUT_1_28(21) => 
        \DATA_OUT_1_28[21]\, DATA_OUT_1_28(20) => 
        \DATA_OUT_1_28[20]\, DATA_OUT_1_28(19) => 
        \DATA_OUT_1_28[19]\, DATA_OUT_1_28(18) => 
        \DATA_OUT_1_28[18]\, DATA_OUT_1_28(17) => 
        \DATA_OUT_1_28[17]\, DATA_OUT_1_28(16) => 
        \DATA_OUT_1_28[16]\, DATA_OUT_1_28(15) => 
        \DATA_OUT_1_28[15]\, DATA_OUT_1_28(14) => 
        \DATA_OUT_1_28[14]\, DATA_OUT_1_28(13) => 
        \DATA_OUT_1_28[13]\, DATA_OUT_1_28(12) => 
        \DATA_OUT_1_28[12]\, DATA_OUT_1_28(11) => 
        \DATA_OUT_1_28[11]\, DATA_OUT_1_28(10) => 
        \DATA_OUT_1_28[10]\, DATA_OUT_1_28(9) => 
        \DATA_OUT_1_28[9]\, DATA_OUT_1_28(8) => 
        \DATA_OUT_1_28[8]\, DATA_OUT_1_28(7) => 
        \DATA_OUT_1_28[7]\, DATA_OUT_1_28(6) => 
        \DATA_OUT_1_28[6]\, DATA_OUT_1_28(5) => 
        \DATA_OUT_1_28[5]\, DATA_OUT_1_28(4) => 
        \DATA_OUT_1_28[4]\, DATA_OUT_1_28(3) => 
        \DATA_OUT_1_28[3]\, DATA_OUT_1_28(2) => 
        \DATA_OUT_1_28[2]\, DATA_OUT_1_28(1) => 
        \DATA_OUT_1_28[1]\, DATA_OUT_1_28(0) => 
        \DATA_OUT_1_28[0]\, DATA_OUT_1_29(25) => 
        \DATA_OUT_1_29[25]\, DATA_OUT_1_29(24) => 
        \DATA_OUT_1_29[24]\, DATA_OUT_1_29(23) => 
        \DATA_OUT_1_29[23]\, DATA_OUT_1_29(22) => 
        \DATA_OUT_1_29[22]\, DATA_OUT_1_29(21) => 
        \DATA_OUT_1_29[21]\, DATA_OUT_1_29(20) => 
        \DATA_OUT_1_29[20]\, DATA_OUT_1_29(19) => 
        \DATA_OUT_1_29[19]\, DATA_OUT_1_29(18) => 
        \DATA_OUT_1_29[18]\, DATA_OUT_1_29(17) => 
        \DATA_OUT_1_29[17]\, DATA_OUT_1_29(16) => 
        \DATA_OUT_1_29[16]\, DATA_OUT_1_29(15) => 
        \DATA_OUT_1_29[15]\, DATA_OUT_1_29(14) => 
        \DATA_OUT_1_29[14]\, DATA_OUT_1_29(13) => 
        \DATA_OUT_1_29[13]\, DATA_OUT_1_29(12) => 
        \DATA_OUT_1_29[12]\, DATA_OUT_1_29(11) => 
        \DATA_OUT_1_29[11]\, DATA_OUT_1_29(10) => 
        \DATA_OUT_1_29[10]\, DATA_OUT_1_29(9) => 
        \DATA_OUT_1_29[9]\, DATA_OUT_1_29(8) => 
        \DATA_OUT_1_29[8]\, DATA_OUT_1_29(7) => 
        \DATA_OUT_1_29[7]\, DATA_OUT_1_29(6) => 
        \DATA_OUT_1_29[6]\, DATA_OUT_1_29(5) => 
        \DATA_OUT_1_29[5]\, DATA_OUT_1_29(4) => 
        \DATA_OUT_1_29[4]\, DATA_OUT_1_29(3) => 
        \DATA_OUT_1_29[3]\, DATA_OUT_1_29(2) => 
        \DATA_OUT_1_29[2]\, DATA_OUT_1_29(1) => 
        \DATA_OUT_1_29[1]\, DATA_OUT_1_29(0) => 
        \DATA_OUT_1_29[0]\, DATA_OUT_1_30(25) => 
        \DATA_OUT_1_30[25]\, DATA_OUT_1_30(24) => 
        \DATA_OUT_1_30[24]\, DATA_OUT_1_30(23) => 
        \DATA_OUT_1_30[23]\, DATA_OUT_1_30(22) => 
        \DATA_OUT_1_30[22]\, DATA_OUT_1_30(21) => 
        \DATA_OUT_1_30[21]\, DATA_OUT_1_30(20) => 
        \DATA_OUT_1_30[20]\, DATA_OUT_1_30(19) => 
        \DATA_OUT_1_30[19]\, DATA_OUT_1_30(18) => 
        \DATA_OUT_1_30[18]\, DATA_OUT_1_30(17) => 
        \DATA_OUT_1_30[17]\, DATA_OUT_1_30(16) => 
        \DATA_OUT_1_30[16]\, DATA_OUT_1_30(15) => 
        \DATA_OUT_1_30[15]\, DATA_OUT_1_30(14) => 
        \DATA_OUT_1_30[14]\, DATA_OUT_1_30(13) => 
        \DATA_OUT_1_30[13]\, DATA_OUT_1_30(12) => 
        \DATA_OUT_1_30[12]\, DATA_OUT_1_30(11) => 
        \DATA_OUT_1_30[11]\, DATA_OUT_1_30(10) => 
        \DATA_OUT_1_30[10]\, DATA_OUT_1_30(9) => 
        \DATA_OUT_1_30[9]\, DATA_OUT_1_30(8) => 
        \DATA_OUT_1_30[8]\, DATA_OUT_1_30(7) => 
        \DATA_OUT_1_30[7]\, DATA_OUT_1_30(6) => 
        \DATA_OUT_1_30[6]\, DATA_OUT_1_30(5) => 
        \DATA_OUT_1_30[5]\, DATA_OUT_1_30(4) => 
        \DATA_OUT_1_30[4]\, DATA_OUT_1_30(3) => 
        \DATA_OUT_1_30[3]\, DATA_OUT_1_30(2) => 
        \DATA_OUT_1_30[2]\, DATA_OUT_1_30(1) => 
        \DATA_OUT_1_30[1]\, DATA_OUT_1_30(0) => 
        \DATA_OUT_1_30[0]\, DATA_OUT_1_31(25) => 
        \DATA_OUT_1_31[25]\, DATA_OUT_1_31(24) => 
        \DATA_OUT_1_31[24]\, DATA_OUT_1_31(23) => 
        \DATA_OUT_1_31[23]\, DATA_OUT_1_31(22) => 
        \DATA_OUT_1_31[22]\, DATA_OUT_1_31(21) => 
        \DATA_OUT_1_31[21]\, DATA_OUT_1_31(20) => 
        \DATA_OUT_1_31[20]\, DATA_OUT_1_31(19) => 
        \DATA_OUT_1_31[19]\, DATA_OUT_1_31(18) => 
        \DATA_OUT_1_31[18]\, DATA_OUT_1_31(17) => 
        \DATA_OUT_1_31[17]\, DATA_OUT_1_31(16) => 
        \DATA_OUT_1_31[16]\, DATA_OUT_1_31(15) => 
        \DATA_OUT_1_31[15]\, DATA_OUT_1_31(14) => 
        \DATA_OUT_1_31[14]\, DATA_OUT_1_31(13) => 
        \DATA_OUT_1_31[13]\, DATA_OUT_1_31(12) => 
        \DATA_OUT_1_31[12]\, DATA_OUT_1_31(11) => 
        \DATA_OUT_1_31[11]\, DATA_OUT_1_31(10) => 
        \DATA_OUT_1_31[10]\, DATA_OUT_1_31(9) => 
        \DATA_OUT_1_31[9]\, DATA_OUT_1_31(8) => 
        \DATA_OUT_1_31[8]\, DATA_OUT_1_31(7) => 
        \DATA_OUT_1_31[7]\, DATA_OUT_1_31(6) => 
        \DATA_OUT_1_31[6]\, DATA_OUT_1_31(5) => 
        \DATA_OUT_1_31[5]\, DATA_OUT_1_31(4) => 
        \DATA_OUT_1_31[4]\, DATA_OUT_1_31(3) => 
        \DATA_OUT_1_31[3]\, DATA_OUT_1_31(2) => 
        \DATA_OUT_1_31[2]\, DATA_OUT_1_31(1) => 
        \DATA_OUT_1_31[1]\, DATA_OUT_1_31(0) => 
        \DATA_OUT_1_31[0]\, DATA_OUT_1_32(25) => 
        \DATA_OUT_1_32[25]\, DATA_OUT_1_32(24) => 
        \DATA_OUT_1_32[24]\, DATA_OUT_1_32(23) => 
        \DATA_OUT_1_32[23]\, DATA_OUT_1_32(22) => 
        \DATA_OUT_1_32[22]\, DATA_OUT_1_32(21) => 
        \DATA_OUT_1_32[21]\, DATA_OUT_1_32(20) => 
        \DATA_OUT_1_32[20]\, DATA_OUT_1_32(19) => 
        \DATA_OUT_1_32[19]\, DATA_OUT_1_32(18) => 
        \DATA_OUT_1_32[18]\, DATA_OUT_1_32(17) => 
        \DATA_OUT_1_32[17]\, DATA_OUT_1_32(16) => 
        \DATA_OUT_1_32[16]\, DATA_OUT_1_32(15) => 
        \DATA_OUT_1_32[15]\, DATA_OUT_1_32(14) => 
        \DATA_OUT_1_32[14]\, DATA_OUT_1_32(13) => 
        \DATA_OUT_1_32[13]\, DATA_OUT_1_32(12) => 
        \DATA_OUT_1_32[12]\, DATA_OUT_1_32(11) => 
        \DATA_OUT_1_32[11]\, DATA_OUT_1_32(10) => 
        \DATA_OUT_1_32[10]\, DATA_OUT_1_32(9) => 
        \DATA_OUT_1_32[9]\, DATA_OUT_1_32(8) => 
        \DATA_OUT_1_32[8]\, DATA_OUT_1_32(7) => 
        \DATA_OUT_1_32[7]\, DATA_OUT_1_32(6) => 
        \DATA_OUT_1_32[6]\, DATA_OUT_1_32(5) => 
        \DATA_OUT_1_32[5]\, DATA_OUT_1_32(4) => 
        \DATA_OUT_1_32[4]\, DATA_OUT_1_32(3) => 
        \DATA_OUT_1_32[3]\, DATA_OUT_1_32(2) => 
        \DATA_OUT_1_32[2]\, DATA_OUT_1_32(1) => 
        \DATA_OUT_1_32[1]\, DATA_OUT_1_32(0) => 
        \DATA_OUT_1_32[0]\, DATA_OUT_1_33(25) => 
        \DATA_OUT_1_33[25]\, DATA_OUT_1_33(24) => 
        \DATA_OUT_1_33[24]\, DATA_OUT_1_33(23) => 
        \DATA_OUT_1_33[23]\, DATA_OUT_1_33(22) => 
        \DATA_OUT_1_33[22]\, DATA_OUT_1_33(21) => 
        \DATA_OUT_1_33[21]\, DATA_OUT_1_33(20) => 
        \DATA_OUT_1_33[20]\, DATA_OUT_1_33(19) => 
        \DATA_OUT_1_33[19]\, DATA_OUT_1_33(18) => 
        \DATA_OUT_1_33[18]\, DATA_OUT_1_33(17) => 
        \DATA_OUT_1_33[17]\, DATA_OUT_1_33(16) => 
        \DATA_OUT_1_33[16]\, DATA_OUT_1_33(15) => 
        \DATA_OUT_1_33[15]\, DATA_OUT_1_33(14) => 
        \DATA_OUT_1_33[14]\, DATA_OUT_1_33(13) => 
        \DATA_OUT_1_33[13]\, DATA_OUT_1_33(12) => 
        \DATA_OUT_1_33[12]\, DATA_OUT_1_33(11) => 
        \DATA_OUT_1_33[11]\, DATA_OUT_1_33(10) => 
        \DATA_OUT_1_33[10]\, DATA_OUT_1_33(9) => 
        \DATA_OUT_1_33[9]\, DATA_OUT_1_33(8) => 
        \DATA_OUT_1_33[8]\, DATA_OUT_1_33(7) => 
        \DATA_OUT_1_33[7]\, DATA_OUT_1_33(6) => 
        \DATA_OUT_1_33[6]\, DATA_OUT_1_33(5) => 
        \DATA_OUT_1_33[5]\, DATA_OUT_1_33(4) => 
        \DATA_OUT_1_33[4]\, DATA_OUT_1_33(3) => 
        \DATA_OUT_1_33[3]\, DATA_OUT_1_33(2) => 
        \DATA_OUT_1_33[2]\, DATA_OUT_1_33(1) => 
        \DATA_OUT_1_33[1]\, DATA_OUT_1_33(0) => 
        \DATA_OUT_1_33[0]\, DATA_OUT_1_34(25) => 
        \DATA_OUT_1_34[25]\, DATA_OUT_1_34(24) => 
        \DATA_OUT_1_34[24]\, DATA_OUT_1_34(23) => 
        \DATA_OUT_1_34[23]\, DATA_OUT_1_34(22) => 
        \DATA_OUT_1_34[22]\, DATA_OUT_1_34(21) => 
        \DATA_OUT_1_34[21]\, DATA_OUT_1_34(20) => 
        \DATA_OUT_1_34[20]\, DATA_OUT_1_34(19) => 
        \DATA_OUT_1_34[19]\, DATA_OUT_1_34(18) => 
        \DATA_OUT_1_34[18]\, DATA_OUT_1_34(17) => 
        \DATA_OUT_1_34[17]\, DATA_OUT_1_34(16) => 
        \DATA_OUT_1_34[16]\, DATA_OUT_1_34(15) => 
        \DATA_OUT_1_34[15]\, DATA_OUT_1_34(14) => 
        \DATA_OUT_1_34[14]\, DATA_OUT_1_34(13) => 
        \DATA_OUT_1_34[13]\, DATA_OUT_1_34(12) => 
        \DATA_OUT_1_34[12]\, DATA_OUT_1_34(11) => 
        \DATA_OUT_1_34[11]\, DATA_OUT_1_34(10) => 
        \DATA_OUT_1_34[10]\, DATA_OUT_1_34(9) => 
        \DATA_OUT_1_34[9]\, DATA_OUT_1_34(8) => 
        \DATA_OUT_1_34[8]\, DATA_OUT_1_34(7) => 
        \DATA_OUT_1_34[7]\, DATA_OUT_1_34(6) => 
        \DATA_OUT_1_34[6]\, DATA_OUT_1_34(5) => 
        \DATA_OUT_1_34[5]\, DATA_OUT_1_34(4) => 
        \DATA_OUT_1_34[4]\, DATA_OUT_1_34(3) => 
        \DATA_OUT_1_34[3]\, DATA_OUT_1_34(2) => 
        \DATA_OUT_1_34[2]\, DATA_OUT_1_34(1) => 
        \DATA_OUT_1_34[1]\, DATA_OUT_1_34(0) => 
        \DATA_OUT_1_34[0]\, DATA_OUT_1_35(25) => 
        \DATA_OUT_1_35[25]\, DATA_OUT_1_35(24) => 
        \DATA_OUT_1_35[24]\, DATA_OUT_1_35(23) => 
        \DATA_OUT_1_35[23]\, DATA_OUT_1_35(22) => 
        \DATA_OUT_1_35[22]\, DATA_OUT_1_35(21) => 
        \DATA_OUT_1_35[21]\, DATA_OUT_1_35(20) => 
        \DATA_OUT_1_35[20]\, DATA_OUT_1_35(19) => 
        \DATA_OUT_1_35[19]\, DATA_OUT_1_35(18) => 
        \DATA_OUT_1_35[18]\, DATA_OUT_1_35(17) => 
        \DATA_OUT_1_35[17]\, DATA_OUT_1_35(16) => 
        \DATA_OUT_1_35[16]\, DATA_OUT_1_35(15) => 
        \DATA_OUT_1_35[15]\, DATA_OUT_1_35(14) => 
        \DATA_OUT_1_35[14]\, DATA_OUT_1_35(13) => 
        \DATA_OUT_1_35[13]\, DATA_OUT_1_35(12) => 
        \DATA_OUT_1_35[12]\, DATA_OUT_1_35(11) => 
        \DATA_OUT_1_35[11]\, DATA_OUT_1_35(10) => 
        \DATA_OUT_1_35[10]\, DATA_OUT_1_35(9) => 
        \DATA_OUT_1_35[9]\, DATA_OUT_1_35(8) => 
        \DATA_OUT_1_35[8]\, DATA_OUT_1_35(7) => 
        \DATA_OUT_1_35[7]\, DATA_OUT_1_35(6) => 
        \DATA_OUT_1_35[6]\, DATA_OUT_1_35(5) => 
        \DATA_OUT_1_35[5]\, DATA_OUT_1_35(4) => 
        \DATA_OUT_1_35[4]\, DATA_OUT_1_35(3) => 
        \DATA_OUT_1_35[3]\, DATA_OUT_1_35(2) => 
        \DATA_OUT_1_35[2]\, DATA_OUT_1_35(1) => 
        \DATA_OUT_1_35[1]\, DATA_OUT_1_35(0) => 
        \DATA_OUT_1_35[0]\, DATA_OUT_1_36(25) => 
        \DATA_OUT_1_36[25]\, DATA_OUT_1_36(24) => 
        \DATA_OUT_1_36[24]\, DATA_OUT_1_36(23) => 
        \DATA_OUT_1_36[23]\, DATA_OUT_1_36(22) => 
        \DATA_OUT_1_36[22]\, DATA_OUT_1_36(21) => 
        \DATA_OUT_1_36[21]\, DATA_OUT_1_36(20) => 
        \DATA_OUT_1_36[20]\, DATA_OUT_1_36(19) => 
        \DATA_OUT_1_36[19]\, DATA_OUT_1_36(18) => 
        \DATA_OUT_1_36[18]\, DATA_OUT_1_36(17) => 
        \DATA_OUT_1_36[17]\, DATA_OUT_1_36(16) => 
        \DATA_OUT_1_36[16]\, DATA_OUT_1_36(15) => 
        \DATA_OUT_1_36[15]\, DATA_OUT_1_36(14) => 
        \DATA_OUT_1_36[14]\, DATA_OUT_1_36(13) => 
        \DATA_OUT_1_36[13]\, DATA_OUT_1_36(12) => 
        \DATA_OUT_1_36[12]\, DATA_OUT_1_36(11) => 
        \DATA_OUT_1_36[11]\, DATA_OUT_1_36(10) => 
        \DATA_OUT_1_36[10]\, DATA_OUT_1_36(9) => 
        \DATA_OUT_1_36[9]\, DATA_OUT_1_36(8) => 
        \DATA_OUT_1_36[8]\, DATA_OUT_1_36(7) => 
        \DATA_OUT_1_36[7]\, DATA_OUT_1_36(6) => 
        \DATA_OUT_1_36[6]\, DATA_OUT_1_36(5) => 
        \DATA_OUT_1_36[5]\, DATA_OUT_1_36(4) => 
        \DATA_OUT_1_36[4]\, DATA_OUT_1_36(3) => 
        \DATA_OUT_1_36[3]\, DATA_OUT_1_36(2) => 
        \DATA_OUT_1_36[2]\, DATA_OUT_1_36(1) => 
        \DATA_OUT_1_36[1]\, DATA_OUT_1_36(0) => 
        \DATA_OUT_1_36[0]\, DATA_OUT_1_37(25) => 
        \DATA_OUT_1_37[25]\, DATA_OUT_1_37(24) => 
        \DATA_OUT_1_37[24]\, DATA_OUT_1_37(23) => 
        \DATA_OUT_1_37[23]\, DATA_OUT_1_37(22) => 
        \DATA_OUT_1_37[22]\, DATA_OUT_1_37(21) => 
        \DATA_OUT_1_37[21]\, DATA_OUT_1_37(20) => 
        \DATA_OUT_1_37[20]\, DATA_OUT_1_37(19) => 
        \DATA_OUT_1_37[19]\, DATA_OUT_1_37(18) => 
        \DATA_OUT_1_37[18]\, DATA_OUT_1_37(17) => 
        \DATA_OUT_1_37[17]\, DATA_OUT_1_37(16) => 
        \DATA_OUT_1_37[16]\, DATA_OUT_1_37(15) => 
        \DATA_OUT_1_37[15]\, DATA_OUT_1_37(14) => 
        \DATA_OUT_1_37[14]\, DATA_OUT_1_37(13) => 
        \DATA_OUT_1_37[13]\, DATA_OUT_1_37(12) => 
        \DATA_OUT_1_37[12]\, DATA_OUT_1_37(11) => 
        \DATA_OUT_1_37[11]\, DATA_OUT_1_37(10) => 
        \DATA_OUT_1_37[10]\, DATA_OUT_1_37(9) => 
        \DATA_OUT_1_37[9]\, DATA_OUT_1_37(8) => 
        \DATA_OUT_1_37[8]\, DATA_OUT_1_37(7) => 
        \DATA_OUT_1_37[7]\, DATA_OUT_1_37(6) => 
        \DATA_OUT_1_37[6]\, DATA_OUT_1_37(5) => 
        \DATA_OUT_1_37[5]\, DATA_OUT_1_37(4) => 
        \DATA_OUT_1_37[4]\, DATA_OUT_1_37(3) => 
        \DATA_OUT_1_37[3]\, DATA_OUT_1_37(2) => 
        \DATA_OUT_1_37[2]\, DATA_OUT_1_37(1) => 
        \DATA_OUT_1_37[1]\, DATA_OUT_1_37(0) => 
        \DATA_OUT_1_37[0]\, DATA_OUT_1_38(25) => 
        \DATA_OUT_1_38[25]\, DATA_OUT_1_38(24) => 
        \DATA_OUT_1_38[24]\, DATA_OUT_1_38(23) => 
        \DATA_OUT_1_38[23]\, DATA_OUT_1_38(22) => 
        \DATA_OUT_1_38[22]\, DATA_OUT_1_38(21) => 
        \DATA_OUT_1_38[21]\, DATA_OUT_1_38(20) => 
        \DATA_OUT_1_38[20]\, DATA_OUT_1_38(19) => 
        \DATA_OUT_1_38[19]\, DATA_OUT_1_38(18) => 
        \DATA_OUT_1_38[18]\, DATA_OUT_1_38(17) => 
        \DATA_OUT_1_38[17]\, DATA_OUT_1_38(16) => 
        \DATA_OUT_1_38[16]\, DATA_OUT_1_38(15) => 
        \DATA_OUT_1_38[15]\, DATA_OUT_1_38(14) => 
        \DATA_OUT_1_38[14]\, DATA_OUT_1_38(13) => 
        \DATA_OUT_1_38[13]\, DATA_OUT_1_38(12) => 
        \DATA_OUT_1_38[12]\, DATA_OUT_1_38(11) => 
        \DATA_OUT_1_38[11]\, DATA_OUT_1_38(10) => 
        \DATA_OUT_1_38[10]\, DATA_OUT_1_38(9) => 
        \DATA_OUT_1_38[9]\, DATA_OUT_1_38(8) => 
        \DATA_OUT_1_38[8]\, DATA_OUT_1_38(7) => 
        \DATA_OUT_1_38[7]\, DATA_OUT_1_38(6) => 
        \DATA_OUT_1_38[6]\, DATA_OUT_1_38(5) => 
        \DATA_OUT_1_38[5]\, DATA_OUT_1_38(4) => 
        \DATA_OUT_1_38[4]\, DATA_OUT_1_38(3) => 
        \DATA_OUT_1_38[3]\, DATA_OUT_1_38(2) => 
        \DATA_OUT_1_38[2]\, DATA_OUT_1_38(1) => 
        \DATA_OUT_1_38[1]\, DATA_OUT_1_38(0) => 
        \DATA_OUT_1_38[0]\, DATA_OUT_1_39(25) => 
        \DATA_OUT_1_39[25]\, DATA_OUT_1_39(24) => 
        \DATA_OUT_1_39[24]\, DATA_OUT_1_39(23) => 
        \DATA_OUT_1_39[23]\, DATA_OUT_1_39(22) => 
        \DATA_OUT_1_39[22]\, DATA_OUT_1_39(21) => 
        \DATA_OUT_1_39[21]\, DATA_OUT_1_39(20) => 
        \DATA_OUT_1_39[20]\, DATA_OUT_1_39(19) => 
        \DATA_OUT_1_39[19]\, DATA_OUT_1_39(18) => 
        \DATA_OUT_1_39[18]\, DATA_OUT_1_39(17) => 
        \DATA_OUT_1_39[17]\, DATA_OUT_1_39(16) => 
        \DATA_OUT_1_39[16]\, DATA_OUT_1_39(15) => 
        \DATA_OUT_1_39[15]\, DATA_OUT_1_39(14) => 
        \DATA_OUT_1_39[14]\, DATA_OUT_1_39(13) => 
        \DATA_OUT_1_39[13]\, DATA_OUT_1_39(12) => 
        \DATA_OUT_1_39[12]\, DATA_OUT_1_39(11) => 
        \DATA_OUT_1_39[11]\, DATA_OUT_1_39(10) => 
        \DATA_OUT_1_39[10]\, DATA_OUT_1_39(9) => 
        \DATA_OUT_1_39[9]\, DATA_OUT_1_39(8) => 
        \DATA_OUT_1_39[8]\, DATA_OUT_1_39(7) => 
        \DATA_OUT_1_39[7]\, DATA_OUT_1_39(6) => 
        \DATA_OUT_1_39[6]\, DATA_OUT_1_39(5) => 
        \DATA_OUT_1_39[5]\, DATA_OUT_1_39(4) => 
        \DATA_OUT_1_39[4]\, DATA_OUT_1_39(3) => 
        \DATA_OUT_1_39[3]\, DATA_OUT_1_39(2) => 
        \DATA_OUT_1_39[2]\, DATA_OUT_1_39(1) => 
        \DATA_OUT_1_39[1]\, DATA_OUT_1_39(0) => 
        \DATA_OUT_1_39[0]\, DATA_OUT_1_40(25) => 
        \DATA_OUT_1_40[25]\, DATA_OUT_1_40(24) => 
        \DATA_OUT_1_40[24]\, DATA_OUT_1_40(23) => 
        \DATA_OUT_1_40[23]\, DATA_OUT_1_40(22) => 
        \DATA_OUT_1_40[22]\, DATA_OUT_1_40(21) => 
        \DATA_OUT_1_40[21]\, DATA_OUT_1_40(20) => 
        \DATA_OUT_1_40[20]\, DATA_OUT_1_40(19) => 
        \DATA_OUT_1_40[19]\, DATA_OUT_1_40(18) => 
        \DATA_OUT_1_40[18]\, DATA_OUT_1_40(17) => 
        \DATA_OUT_1_40[17]\, DATA_OUT_1_40(16) => 
        \DATA_OUT_1_40[16]\, DATA_OUT_1_40(15) => 
        \DATA_OUT_1_40[15]\, DATA_OUT_1_40(14) => 
        \DATA_OUT_1_40[14]\, DATA_OUT_1_40(13) => 
        \DATA_OUT_1_40[13]\, DATA_OUT_1_40(12) => 
        \DATA_OUT_1_40[12]\, DATA_OUT_1_40(11) => 
        \DATA_OUT_1_40[11]\, DATA_OUT_1_40(10) => 
        \DATA_OUT_1_40[10]\, DATA_OUT_1_40(9) => 
        \DATA_OUT_1_40[9]\, DATA_OUT_1_40(8) => 
        \DATA_OUT_1_40[8]\, DATA_OUT_1_40(7) => 
        \DATA_OUT_1_40[7]\, DATA_OUT_1_40(6) => 
        \DATA_OUT_1_40[6]\, DATA_OUT_1_40(5) => 
        \DATA_OUT_1_40[5]\, DATA_OUT_1_40(4) => 
        \DATA_OUT_1_40[4]\, DATA_OUT_1_40(3) => 
        \DATA_OUT_1_40[3]\, DATA_OUT_1_40(2) => 
        \DATA_OUT_1_40[2]\, DATA_OUT_1_40(1) => 
        \DATA_OUT_1_40[1]\, DATA_OUT_1_40(0) => 
        \DATA_OUT_1_40[0]\, DATA_OUT_1_41(25) => 
        \DATA_OUT_1_41[25]\, DATA_OUT_1_41(24) => 
        \DATA_OUT_1_41[24]\, DATA_OUT_1_41(23) => 
        \DATA_OUT_1_41[23]\, DATA_OUT_1_41(22) => 
        \DATA_OUT_1_41[22]\, DATA_OUT_1_41(21) => 
        \DATA_OUT_1_41[21]\, DATA_OUT_1_41(20) => 
        \DATA_OUT_1_41[20]\, DATA_OUT_1_41(19) => 
        \DATA_OUT_1_41[19]\, DATA_OUT_1_41(18) => 
        \DATA_OUT_1_41[18]\, DATA_OUT_1_41(17) => 
        \DATA_OUT_1_41[17]\, DATA_OUT_1_41(16) => 
        \DATA_OUT_1_41[16]\, DATA_OUT_1_41(15) => 
        \DATA_OUT_1_41[15]\, DATA_OUT_1_41(14) => 
        \DATA_OUT_1_41[14]\, DATA_OUT_1_41(13) => 
        \DATA_OUT_1_41[13]\, DATA_OUT_1_41(12) => 
        \DATA_OUT_1_41[12]\, DATA_OUT_1_41(11) => 
        \DATA_OUT_1_41[11]\, DATA_OUT_1_41(10) => 
        \DATA_OUT_1_41[10]\, DATA_OUT_1_41(9) => 
        \DATA_OUT_1_41[9]\, DATA_OUT_1_41(8) => 
        \DATA_OUT_1_41[8]\, DATA_OUT_1_41(7) => 
        \DATA_OUT_1_41[7]\, DATA_OUT_1_41(6) => 
        \DATA_OUT_1_41[6]\, DATA_OUT_1_41(5) => 
        \DATA_OUT_1_41[5]\, DATA_OUT_1_41(4) => 
        \DATA_OUT_1_41[4]\, DATA_OUT_1_41(3) => 
        \DATA_OUT_1_41[3]\, DATA_OUT_1_41(2) => 
        \DATA_OUT_1_41[2]\, DATA_OUT_1_41(1) => 
        \DATA_OUT_1_41[1]\, DATA_OUT_1_41(0) => 
        \DATA_OUT_1_41[0]\, DATA_OUT_1_42(25) => 
        \DATA_OUT_1_42[25]\, DATA_OUT_1_42(24) => 
        \DATA_OUT_1_42[24]\, DATA_OUT_1_42(23) => 
        \DATA_OUT_1_42[23]\, DATA_OUT_1_42(22) => 
        \DATA_OUT_1_42[22]\, DATA_OUT_1_42(21) => 
        \DATA_OUT_1_42[21]\, DATA_OUT_1_42(20) => 
        \DATA_OUT_1_42[20]\, DATA_OUT_1_42(19) => 
        \DATA_OUT_1_42[19]\, DATA_OUT_1_42(18) => 
        \DATA_OUT_1_42[18]\, DATA_OUT_1_42(17) => 
        \DATA_OUT_1_42[17]\, DATA_OUT_1_42(16) => 
        \DATA_OUT_1_42[16]\, DATA_OUT_1_42(15) => 
        \DATA_OUT_1_42[15]\, DATA_OUT_1_42(14) => 
        \DATA_OUT_1_42[14]\, DATA_OUT_1_42(13) => 
        \DATA_OUT_1_42[13]\, DATA_OUT_1_42(12) => 
        \DATA_OUT_1_42[12]\, DATA_OUT_1_42(11) => 
        \DATA_OUT_1_42[11]\, DATA_OUT_1_42(10) => 
        \DATA_OUT_1_42[10]\, DATA_OUT_1_42(9) => 
        \DATA_OUT_1_42[9]\, DATA_OUT_1_42(8) => 
        \DATA_OUT_1_42[8]\, DATA_OUT_1_42(7) => 
        \DATA_OUT_1_42[7]\, DATA_OUT_1_42(6) => 
        \DATA_OUT_1_42[6]\, DATA_OUT_1_42(5) => 
        \DATA_OUT_1_42[5]\, DATA_OUT_1_42(4) => 
        \DATA_OUT_1_42[4]\, DATA_OUT_1_42(3) => 
        \DATA_OUT_1_42[3]\, DATA_OUT_1_42(2) => 
        \DATA_OUT_1_42[2]\, DATA_OUT_1_42(1) => 
        \DATA_OUT_1_42[1]\, DATA_OUT_1_42(0) => 
        \DATA_OUT_1_42[0]\, DATA_OUT_1_43(25) => 
        \DATA_OUT_1_43[25]\, DATA_OUT_1_43(24) => 
        \DATA_OUT_1_43[24]\, DATA_OUT_1_43(23) => 
        \DATA_OUT_1_43[23]\, DATA_OUT_1_43(22) => 
        \DATA_OUT_1_43[22]\, DATA_OUT_1_43(21) => 
        \DATA_OUT_1_43[21]\, DATA_OUT_1_43(20) => 
        \DATA_OUT_1_43[20]\, DATA_OUT_1_43(19) => 
        \DATA_OUT_1_43[19]\, DATA_OUT_1_43(18) => 
        \DATA_OUT_1_43[18]\, DATA_OUT_1_43(17) => 
        \DATA_OUT_1_43[17]\, DATA_OUT_1_43(16) => 
        \DATA_OUT_1_43[16]\, DATA_OUT_1_43(15) => 
        \DATA_OUT_1_43[15]\, DATA_OUT_1_43(14) => 
        \DATA_OUT_1_43[14]\, DATA_OUT_1_43(13) => 
        \DATA_OUT_1_43[13]\, DATA_OUT_1_43(12) => 
        \DATA_OUT_1_43[12]\, DATA_OUT_1_43(11) => 
        \DATA_OUT_1_43[11]\, DATA_OUT_1_43(10) => 
        \DATA_OUT_1_43[10]\, DATA_OUT_1_43(9) => 
        \DATA_OUT_1_43[9]\, DATA_OUT_1_43(8) => 
        \DATA_OUT_1_43[8]\, DATA_OUT_1_43(7) => 
        \DATA_OUT_1_43[7]\, DATA_OUT_1_43(6) => 
        \DATA_OUT_1_43[6]\, DATA_OUT_1_43(5) => 
        \DATA_OUT_1_43[5]\, DATA_OUT_1_43(4) => 
        \DATA_OUT_1_43[4]\, DATA_OUT_1_43(3) => 
        \DATA_OUT_1_43[3]\, DATA_OUT_1_43(2) => 
        \DATA_OUT_1_43[2]\, DATA_OUT_1_43(1) => 
        \DATA_OUT_1_43[1]\, DATA_OUT_1_43(0) => 
        \DATA_OUT_1_43[0]\, DATA_OUT_1_44(25) => 
        \DATA_OUT_1_44[25]\, DATA_OUT_1_44(24) => 
        \DATA_OUT_1_44[24]\, DATA_OUT_1_44(23) => 
        \DATA_OUT_1_44[23]\, DATA_OUT_1_44(22) => 
        \DATA_OUT_1_44[22]\, DATA_OUT_1_44(21) => 
        \DATA_OUT_1_44[21]\, DATA_OUT_1_44(20) => 
        \DATA_OUT_1_44[20]\, DATA_OUT_1_44(19) => 
        \DATA_OUT_1_44[19]\, DATA_OUT_1_44(18) => 
        \DATA_OUT_1_44[18]\, DATA_OUT_1_44(17) => 
        \DATA_OUT_1_44[17]\, DATA_OUT_1_44(16) => 
        \DATA_OUT_1_44[16]\, DATA_OUT_1_44(15) => 
        \DATA_OUT_1_44[15]\, DATA_OUT_1_44(14) => 
        \DATA_OUT_1_44[14]\, DATA_OUT_1_44(13) => 
        \DATA_OUT_1_44[13]\, DATA_OUT_1_44(12) => 
        \DATA_OUT_1_44[12]\, DATA_OUT_1_44(11) => 
        \DATA_OUT_1_44[11]\, DATA_OUT_1_44(10) => 
        \DATA_OUT_1_44[10]\, DATA_OUT_1_44(9) => 
        \DATA_OUT_1_44[9]\, DATA_OUT_1_44(8) => 
        \DATA_OUT_1_44[8]\, DATA_OUT_1_44(7) => 
        \DATA_OUT_1_44[7]\, DATA_OUT_1_44(6) => 
        \DATA_OUT_1_44[6]\, DATA_OUT_1_44(5) => 
        \DATA_OUT_1_44[5]\, DATA_OUT_1_44(4) => 
        \DATA_OUT_1_44[4]\, DATA_OUT_1_44(3) => 
        \DATA_OUT_1_44[3]\, DATA_OUT_1_44(2) => 
        \DATA_OUT_1_44[2]\, DATA_OUT_1_44(1) => 
        \DATA_OUT_1_44[1]\, DATA_OUT_1_44(0) => 
        \DATA_OUT_1_44[0]\, DATA_OUT_1_45(25) => 
        \DATA_OUT_1_45[25]\, DATA_OUT_1_45(24) => 
        \DATA_OUT_1_45[24]\, DATA_OUT_1_45(23) => 
        \DATA_OUT_1_45[23]\, DATA_OUT_1_45(22) => 
        \DATA_OUT_1_45[22]\, DATA_OUT_1_45(21) => 
        \DATA_OUT_1_45[21]\, DATA_OUT_1_45(20) => 
        \DATA_OUT_1_45[20]\, DATA_OUT_1_45(19) => 
        \DATA_OUT_1_45[19]\, DATA_OUT_1_45(18) => 
        \DATA_OUT_1_45[18]\, DATA_OUT_1_45(17) => 
        \DATA_OUT_1_45[17]\, DATA_OUT_1_45(16) => 
        \DATA_OUT_1_45[16]\, DATA_OUT_1_45(15) => 
        \DATA_OUT_1_45[15]\, DATA_OUT_1_45(14) => 
        \DATA_OUT_1_45[14]\, DATA_OUT_1_45(13) => 
        \DATA_OUT_1_45[13]\, DATA_OUT_1_45(12) => 
        \DATA_OUT_1_45[12]\, DATA_OUT_1_45(11) => 
        \DATA_OUT_1_45[11]\, DATA_OUT_1_45(10) => 
        \DATA_OUT_1_45[10]\, DATA_OUT_1_45(9) => 
        \DATA_OUT_1_45[9]\, DATA_OUT_1_45(8) => 
        \DATA_OUT_1_45[8]\, DATA_OUT_1_45(7) => 
        \DATA_OUT_1_45[7]\, DATA_OUT_1_45(6) => 
        \DATA_OUT_1_45[6]\, DATA_OUT_1_45(5) => 
        \DATA_OUT_1_45[5]\, DATA_OUT_1_45(4) => 
        \DATA_OUT_1_45[4]\, DATA_OUT_1_45(3) => 
        \DATA_OUT_1_45[3]\, DATA_OUT_1_45(2) => 
        \DATA_OUT_1_45[2]\, DATA_OUT_1_45(1) => 
        \DATA_OUT_1_45[1]\, DATA_OUT_1_45(0) => 
        \DATA_OUT_1_45[0]\, DATA_OUT_1_46(25) => 
        \DATA_OUT_1_46[25]\, DATA_OUT_1_46(24) => 
        \DATA_OUT_1_46[24]\, DATA_OUT_1_46(23) => 
        \DATA_OUT_1_46[23]\, DATA_OUT_1_46(22) => 
        \DATA_OUT_1_46[22]\, DATA_OUT_1_46(21) => 
        \DATA_OUT_1_46[21]\, DATA_OUT_1_46(20) => 
        \DATA_OUT_1_46[20]\, DATA_OUT_1_46(19) => 
        \DATA_OUT_1_46[19]\, DATA_OUT_1_46(18) => 
        \DATA_OUT_1_46[18]\, DATA_OUT_1_46(17) => 
        \DATA_OUT_1_46[17]\, DATA_OUT_1_46(16) => 
        \DATA_OUT_1_46[16]\, DATA_OUT_1_46(15) => 
        \DATA_OUT_1_46[15]\, DATA_OUT_1_46(14) => 
        \DATA_OUT_1_46[14]\, DATA_OUT_1_46(13) => 
        \DATA_OUT_1_46[13]\, DATA_OUT_1_46(12) => 
        \DATA_OUT_1_46[12]\, DATA_OUT_1_46(11) => 
        \DATA_OUT_1_46[11]\, DATA_OUT_1_46(10) => 
        \DATA_OUT_1_46[10]\, DATA_OUT_1_46(9) => 
        \DATA_OUT_1_46[9]\, DATA_OUT_1_46(8) => 
        \DATA_OUT_1_46[8]\, DATA_OUT_1_46(7) => 
        \DATA_OUT_1_46[7]\, DATA_OUT_1_46(6) => 
        \DATA_OUT_1_46[6]\, DATA_OUT_1_46(5) => 
        \DATA_OUT_1_46[5]\, DATA_OUT_1_46(4) => 
        \DATA_OUT_1_46[4]\, DATA_OUT_1_46(3) => 
        \DATA_OUT_1_46[3]\, DATA_OUT_1_46(2) => 
        \DATA_OUT_1_46[2]\, DATA_OUT_1_46(1) => 
        \DATA_OUT_1_46[1]\, DATA_OUT_1_46(0) => 
        \DATA_OUT_1_46[0]\, DATA_OUT_1_47(25) => 
        \DATA_OUT_1_47[25]\, DATA_OUT_1_47(24) => 
        \DATA_OUT_1_47[24]\, DATA_OUT_1_47(23) => 
        \DATA_OUT_1_47[23]\, DATA_OUT_1_47(22) => 
        \DATA_OUT_1_47[22]\, DATA_OUT_1_47(21) => 
        \DATA_OUT_1_47[21]\, DATA_OUT_1_47(20) => 
        \DATA_OUT_1_47[20]\, DATA_OUT_1_47(19) => 
        \DATA_OUT_1_47[19]\, DATA_OUT_1_47(18) => 
        \DATA_OUT_1_47[18]\, DATA_OUT_1_47(17) => 
        \DATA_OUT_1_47[17]\, DATA_OUT_1_47(16) => 
        \DATA_OUT_1_47[16]\, DATA_OUT_1_47(15) => 
        \DATA_OUT_1_47[15]\, DATA_OUT_1_47(14) => 
        \DATA_OUT_1_47[14]\, DATA_OUT_1_47(13) => 
        \DATA_OUT_1_47[13]\, DATA_OUT_1_47(12) => 
        \DATA_OUT_1_47[12]\, DATA_OUT_1_47(11) => 
        \DATA_OUT_1_47[11]\, DATA_OUT_1_47(10) => 
        \DATA_OUT_1_47[10]\, DATA_OUT_1_47(9) => 
        \DATA_OUT_1_47[9]\, DATA_OUT_1_47(8) => 
        \DATA_OUT_1_47[8]\, DATA_OUT_1_47(7) => 
        \DATA_OUT_1_47[7]\, DATA_OUT_1_47(6) => 
        \DATA_OUT_1_47[6]\, DATA_OUT_1_47(5) => 
        \DATA_OUT_1_47[5]\, DATA_OUT_1_47(4) => 
        \DATA_OUT_1_47[4]\, DATA_OUT_1_47(3) => 
        \DATA_OUT_1_47[3]\, DATA_OUT_1_47(2) => 
        \DATA_OUT_1_47[2]\, DATA_OUT_1_47(1) => 
        \DATA_OUT_1_47[1]\, DATA_OUT_1_47(0) => 
        \DATA_OUT_1_47[0]\, DATA_OUT_1_48(25) => 
        \DATA_OUT_1_48[25]\, DATA_OUT_1_48(24) => 
        \DATA_OUT_1_48[24]\, DATA_OUT_1_48(23) => 
        \DATA_OUT_1_48[23]\, DATA_OUT_1_48(22) => 
        \DATA_OUT_1_48[22]\, DATA_OUT_1_48(21) => 
        \DATA_OUT_1_48[21]\, DATA_OUT_1_48(20) => 
        \DATA_OUT_1_48[20]\, DATA_OUT_1_48(19) => 
        \DATA_OUT_1_48[19]\, DATA_OUT_1_48(18) => 
        \DATA_OUT_1_48[18]\, DATA_OUT_1_48(17) => 
        \DATA_OUT_1_48[17]\, DATA_OUT_1_48(16) => 
        \DATA_OUT_1_48[16]\, DATA_OUT_1_48(15) => 
        \DATA_OUT_1_48[15]\, DATA_OUT_1_48(14) => 
        \DATA_OUT_1_48[14]\, DATA_OUT_1_48(13) => 
        \DATA_OUT_1_48[13]\, DATA_OUT_1_48(12) => 
        \DATA_OUT_1_48[12]\, DATA_OUT_1_48(11) => 
        \DATA_OUT_1_48[11]\, DATA_OUT_1_48(10) => 
        \DATA_OUT_1_48[10]\, DATA_OUT_1_48(9) => 
        \DATA_OUT_1_48[9]\, DATA_OUT_1_48(8) => 
        \DATA_OUT_1_48[8]\, DATA_OUT_1_48(7) => 
        \DATA_OUT_1_48[7]\, DATA_OUT_1_48(6) => 
        \DATA_OUT_1_48[6]\, DATA_OUT_1_48(5) => 
        \DATA_OUT_1_48[5]\, DATA_OUT_1_48(4) => 
        \DATA_OUT_1_48[4]\, DATA_OUT_1_48(3) => 
        \DATA_OUT_1_48[3]\, DATA_OUT_1_48(2) => 
        \DATA_OUT_1_48[2]\, DATA_OUT_1_48(1) => 
        \DATA_OUT_1_48[1]\, DATA_OUT_1_48(0) => 
        \DATA_OUT_1_48[0]\, DATA_OUT_1_49(25) => 
        \DATA_OUT_1_49[25]\, DATA_OUT_1_49(24) => 
        \DATA_OUT_1_49[24]\, DATA_OUT_1_49(23) => 
        \DATA_OUT_1_49[23]\, DATA_OUT_1_49(22) => 
        \DATA_OUT_1_49[22]\, DATA_OUT_1_49(21) => 
        \DATA_OUT_1_49[21]\, DATA_OUT_1_49(20) => 
        \DATA_OUT_1_49[20]\, DATA_OUT_1_49(19) => 
        \DATA_OUT_1_49[19]\, DATA_OUT_1_49(18) => 
        \DATA_OUT_1_49[18]\, DATA_OUT_1_49(17) => 
        \DATA_OUT_1_49[17]\, DATA_OUT_1_49(16) => 
        \DATA_OUT_1_49[16]\, DATA_OUT_1_49(15) => 
        \DATA_OUT_1_49[15]\, DATA_OUT_1_49(14) => 
        \DATA_OUT_1_49[14]\, DATA_OUT_1_49(13) => 
        \DATA_OUT_1_49[13]\, DATA_OUT_1_49(12) => 
        \DATA_OUT_1_49[12]\, DATA_OUT_1_49(11) => 
        \DATA_OUT_1_49[11]\, DATA_OUT_1_49(10) => 
        \DATA_OUT_1_49[10]\, DATA_OUT_1_49(9) => 
        \DATA_OUT_1_49[9]\, DATA_OUT_1_49(8) => 
        \DATA_OUT_1_49[8]\, DATA_OUT_1_49(7) => 
        \DATA_OUT_1_49[7]\, DATA_OUT_1_49(6) => 
        \DATA_OUT_1_49[6]\, DATA_OUT_1_49(5) => 
        \DATA_OUT_1_49[5]\, DATA_OUT_1_49(4) => 
        \DATA_OUT_1_49[4]\, DATA_OUT_1_49(3) => 
        \DATA_OUT_1_49[3]\, DATA_OUT_1_49(2) => 
        \DATA_OUT_1_49[2]\, DATA_OUT_1_49(1) => 
        \DATA_OUT_1_49[1]\, DATA_OUT_1_49(0) => 
        \DATA_OUT_1_49[0]\, DATA_OUT_1_50(25) => 
        \DATA_OUT_1_50[25]\, DATA_OUT_1_50(24) => 
        \DATA_OUT_1_50[24]\, DATA_OUT_1_50(23) => 
        \DATA_OUT_1_50[23]\, DATA_OUT_1_50(22) => 
        \DATA_OUT_1_50[22]\, DATA_OUT_1_50(21) => 
        \DATA_OUT_1_50[21]\, DATA_OUT_1_50(20) => 
        \DATA_OUT_1_50[20]\, DATA_OUT_1_50(19) => 
        \DATA_OUT_1_50[19]\, DATA_OUT_1_50(18) => 
        \DATA_OUT_1_50[18]\, DATA_OUT_1_50(17) => 
        \DATA_OUT_1_50[17]\, DATA_OUT_1_50(16) => 
        \DATA_OUT_1_50[16]\, DATA_OUT_1_50(15) => 
        \DATA_OUT_1_50[15]\, DATA_OUT_1_50(14) => 
        \DATA_OUT_1_50[14]\, DATA_OUT_1_50(13) => 
        \DATA_OUT_1_50[13]\, DATA_OUT_1_50(12) => 
        \DATA_OUT_1_50[12]\, DATA_OUT_1_50(11) => 
        \DATA_OUT_1_50[11]\, DATA_OUT_1_50(10) => 
        \DATA_OUT_1_50[10]\, DATA_OUT_1_50(9) => 
        \DATA_OUT_1_50[9]\, DATA_OUT_1_50(8) => 
        \DATA_OUT_1_50[8]\, DATA_OUT_1_50(7) => 
        \DATA_OUT_1_50[7]\, DATA_OUT_1_50(6) => 
        \DATA_OUT_1_50[6]\, DATA_OUT_1_50(5) => 
        \DATA_OUT_1_50[5]\, DATA_OUT_1_50(4) => 
        \DATA_OUT_1_50[4]\, DATA_OUT_1_50(3) => 
        \DATA_OUT_1_50[3]\, DATA_OUT_1_50(2) => 
        \DATA_OUT_1_50[2]\, DATA_OUT_1_50(1) => 
        \DATA_OUT_1_50[1]\, DATA_OUT_1_50(0) => 
        \DATA_OUT_1_50[0]\, DATA_OUT_1_51(25) => 
        \DATA_OUT_1_51[25]\, DATA_OUT_1_51(24) => 
        \DATA_OUT_1_51[24]\, DATA_OUT_1_51(23) => 
        \DATA_OUT_1_51[23]\, DATA_OUT_1_51(22) => 
        \DATA_OUT_1_51[22]\, DATA_OUT_1_51(21) => 
        \DATA_OUT_1_51[21]\, DATA_OUT_1_51(20) => 
        \DATA_OUT_1_51[20]\, DATA_OUT_1_51(19) => 
        \DATA_OUT_1_51[19]\, DATA_OUT_1_51(18) => 
        \DATA_OUT_1_51[18]\, DATA_OUT_1_51(17) => 
        \DATA_OUT_1_51[17]\, DATA_OUT_1_51(16) => 
        \DATA_OUT_1_51[16]\, DATA_OUT_1_51(15) => 
        \DATA_OUT_1_51[15]\, DATA_OUT_1_51(14) => 
        \DATA_OUT_1_51[14]\, DATA_OUT_1_51(13) => 
        \DATA_OUT_1_51[13]\, DATA_OUT_1_51(12) => 
        \DATA_OUT_1_51[12]\, DATA_OUT_1_51(11) => 
        \DATA_OUT_1_51[11]\, DATA_OUT_1_51(10) => 
        \DATA_OUT_1_51[10]\, DATA_OUT_1_51(9) => 
        \DATA_OUT_1_51[9]\, DATA_OUT_1_51(8) => 
        \DATA_OUT_1_51[8]\, DATA_OUT_1_51(7) => 
        \DATA_OUT_1_51[7]\, DATA_OUT_1_51(6) => 
        \DATA_OUT_1_51[6]\, DATA_OUT_1_51(5) => 
        \DATA_OUT_1_51[5]\, DATA_OUT_1_51(4) => 
        \DATA_OUT_1_51[4]\, DATA_OUT_1_51(3) => 
        \DATA_OUT_1_51[3]\, DATA_OUT_1_51(2) => 
        \DATA_OUT_1_51[2]\, DATA_OUT_1_51(1) => 
        \DATA_OUT_1_51[1]\, DATA_OUT_1_51(0) => 
        \DATA_OUT_1_51[0]\);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 
